`timescale 1 ns/100 ps
// Version: v11.6 SP1 11.6.1.6


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module COREAPB3_MUXPTOB3(
       CoreAPB3_0_APBmslave2_PRDATA,
       CoreAPB3_0_APBmslave3_PRDATA,
       iPSELS_0,
       iPSELS_0_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_1,
       CoreAPB3_0_APBmslave0_PRDATA_m_2,
       CoreAPB3_0_APBmslave1_PRDATA_m,
       CoreAPB3_0_APBmslave4_PRDATA,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       sercon_0,
       sercon_2,
       CoreAPB3_0_APBmslave0_PADDR_0,
       CoreAPB3_0_APBmslave0_PADDR_7,
       serdat_0,
       serdat_2,
       CoreAPB3_0_APBmslave0_PRDATA_m_0_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_4,
       CoreAPB3_0_APBmslave0_PRDATA_m_5,
       CoreAPB3_0_APBmslave0_PRDATA_m_3,
       CoreAPB3_0_APBmslave0_PRDATA_m_2_d0,
       un4_PRDATA_1,
       controlReg14_3,
       CoreAPB3_0_APBmslave0_PSELx,
       r_N_4_mux,
       un12_PSELi,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_0_APBmslave2_PSELx,
       un4_PRDATA,
       un1_PRDATA,
       PRDATA_regif_sn_N_39_mux,
       un14_PRDATA,
       PRDATA_regif_sn_N_26,
       N_809,
       N_829,
       N_810,
       N_830,
       N_807,
       N_827,
       N_808,
       N_828,
       N_812,
       N_832,
       N_806,
       N_826,
       N_813,
       N_833,
       N_811,
       N_831,
       N_840,
       N_842,
       N_837,
       N_841,
       N_839,
       N_838
    );
input  [7:0] CoreAPB3_0_APBmslave2_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [4:4] iPSELS_0;
input  [4:4] iPSELS_0_0;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_0;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_1;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_2;
input  [1:0] CoreAPB3_0_APBmslave1_PRDATA_m;
input  [1:0] CoreAPB3_0_APBmslave4_PRDATA;
output [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
input  sercon_0;
input  sercon_2;
input  CoreAPB3_0_APBmslave0_PADDR_0;
input  CoreAPB3_0_APBmslave0_PADDR_7;
input  serdat_0;
input  serdat_2;
input  CoreAPB3_0_APBmslave0_PRDATA_m_0_d0;
input  CoreAPB3_0_APBmslave0_PRDATA_m_4;
input  CoreAPB3_0_APBmslave0_PRDATA_m_5;
input  CoreAPB3_0_APBmslave0_PRDATA_m_3;
input  CoreAPB3_0_APBmslave0_PRDATA_m_2_d0;
input  un4_PRDATA_1;
input  controlReg14_3;
input  CoreAPB3_0_APBmslave0_PSELx;
output r_N_4_mux;
input  un12_PSELi;
input  CoreAPB3_0_APBmslave3_PSELx;
input  CoreAPB3_0_APBmslave2_PSELx;
input  un4_PRDATA;
input  un1_PRDATA;
input  PRDATA_regif_sn_N_39_mux;
input  un14_PRDATA;
input  PRDATA_regif_sn_N_26;
input  N_809;
input  N_829;
input  N_810;
input  N_830;
input  N_807;
input  N_827;
input  N_808;
input  N_828;
input  N_812;
input  N_832;
input  N_806;
input  N_826;
input  N_813;
input  N_833;
input  N_811;
input  N_831;
input  N_840;
input  N_842;
input  N_837;
input  N_841;
input  N_839;
input  N_838;

    wire PRDATA_m3_0_0_net_1, \PRDATA_0_iv_0[1]_net_1 , 
        \PRDATA_0_iv_0[0]_net_1 , \PRDATA_0_iv_0[2]_net_1 , 
        \PRDATA_0_iv_0[7]_net_1 , \PRDATA_0_iv_0[3]_net_1 , 
        \PRDATA_0_iv_0[6]_net_1 , \PRDATA_0_iv_0[5]_net_1 , 
        \PRDATA_0_iv_0[4]_net_1 , \PRDATA_0_iv_2_a1[0]_net_1 , 
        \PRDATA_0_iv_2_a0[0]_net_1 , \PRDATA_0_iv_1[2]_net_1 , 
        \PRDATA_0[8] , PRDATA_m3_0_d_net_1, \PRDATA_0_iv_1[7]_net_1 , 
        \PRDATA_0_iv_2[1]_net_1 , \PRDATA_0_iv_3[0]_net_1 , GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[1]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[1]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[1]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[1]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \PRDATA_0[10]  (.A(iPSELS_0[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR_7), .C(PRDATA_regif_sn_N_39_mux), 
        .D(iPSELS_0_0[4]), .Y(\PRDATA_0[8] ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[14]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_812), .C(\PRDATA_0[8] ), .D(N_832), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]));
    CFG4 #( .INIT(16'hFFFE) )  \PRDATA_0_iv_3[0]  (.A(
        CoreAPB3_0_APBmslave1_PRDATA_m[0]), .B(
        \PRDATA_0_iv_0[0]_net_1 ), .C(\PRDATA_0_iv_2_a1[0]_net_1 ), .D(
        \PRDATA_0_iv_2_a0[0]_net_1 ), .Y(\PRDATA_0_iv_3[0]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_1[7]  (.A(
        CoreAPB3_0_APBmslave0_PRDATA_m_0[7]), .B(
        CoreAPB3_0_APBmslave0_PRDATA_m_1[7]), .C(
        \PRDATA_0_iv_0[7]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]), .Y(
        \PRDATA_0_iv_1[7]_net_1 ));
    CFG2 #( .INIT(4'h7) )  PRDATA_m3_0_0 (.A(
        CoreAPB3_0_APBmslave0_PSELx), .B(un12_PSELi), .Y(
        PRDATA_m3_0_0_net_1));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[10]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_808), .C(\PRDATA_0[8] ), .D(N_828), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv[0]  (.A(iPSELS_0_0[4]), .B(
        iPSELS_0[4]), .C(\PRDATA_0_iv_3[0]_net_1 ), .D(
        CoreAPB3_0_APBmslave4_PRDATA[0]), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[8]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_806), .C(\PRDATA_0[8] ), .D(N_826), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]));
    CFG4 #( .INIT(16'hFEEE) )  \PRDATA_0_iv[2]  (.A(
        PRDATA_m3_0_d_net_1), .B(\PRDATA_0_iv_1[2]_net_1 ), .C(
        \PRDATA_0[8] ), .D(N_837), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2]));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[12]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_810), .C(\PRDATA_0[8] ), .D(N_830), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]));
    CFG4 #( .INIT(16'hFFEA) )  \PRDATA_0_iv[3]  (.A(
        \PRDATA_0_iv_0[3]_net_1 ), .B(\PRDATA_0[8] ), .C(N_838), .D(
        CoreAPB3_0_APBmslave0_PRDATA_m_2_d0), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3]));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_0_iv_2_a1_1[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR_0), .B(un4_PRDATA_1), .C(
        controlReg14_3), .D(CoreAPB3_0_APBmslave0_PSELx), .Y(r_N_4_mux)
        );
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[7]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[7]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[7]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[7]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv[5]  (.A(\PRDATA_0[8] ), .B(
        N_840), .C(CoreAPB3_0_APBmslave0_PRDATA_m_4), .D(
        \PRDATA_0_iv_0[5]_net_1 ), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5]));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[0]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[0]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[0]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h00EC) )  PRDATA_m3_0_d (.A(serdat_2), .B(
        un14_PRDATA), .C(un4_PRDATA), .D(PRDATA_m3_0_0_net_1), .Y(
        PRDATA_m3_0_d_net_1));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv_1[2]  (.A(un1_PRDATA), .B(
        sercon_2), .C(\PRDATA_0_iv_0[2]_net_1 ), .D(
        PRDATA_m3_0_0_net_1), .Y(\PRDATA_0_iv_1[2]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[6]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[6]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[6]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[6]_net_1 ));
    CFG4 #( .INIT(16'hFFEA) )  \PRDATA_0_iv[4]  (.A(
        \PRDATA_0_iv_0[4]_net_1 ), .B(\PRDATA_0[8] ), .C(N_839), .D(
        CoreAPB3_0_APBmslave0_PRDATA_m_3), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4]));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[15]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_813), .C(\PRDATA_0[8] ), .D(N_833), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv[1]  (.A(iPSELS_0[4]), .B(
        iPSELS_0_0[4]), .C(\PRDATA_0_iv_2[1]_net_1 ), .D(
        CoreAPB3_0_APBmslave4_PRDATA[1]), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1]));
    CFG4 #( .INIT(16'hFFEA) )  \PRDATA_0_iv[6]  (.A(
        \PRDATA_0_iv_0[6]_net_1 ), .B(\PRDATA_0[8] ), .C(N_841), .D(
        CoreAPB3_0_APBmslave0_PRDATA_m_5), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6]));
    CFG3 #( .INIT(8'hEA) )  \PRDATA_0_iv[7]  (.A(
        \PRDATA_0_iv_1[7]_net_1 ), .B(\PRDATA_0[8] ), .C(N_842), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7]));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[3]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[3]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[3]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[3]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \PRDATA_0_iv_2[1]  (.A(
        CoreAPB3_0_APBmslave1_PRDATA_m[1]), .B(
        \PRDATA_0_iv_0[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PRDATA_m_0_d0), .Y(
        \PRDATA_0_iv_2[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_2_a0[0]  (.A(sercon_0), .B(
        un12_PSELi), .C(un1_PRDATA), .D(CoreAPB3_0_APBmslave0_PSELx), 
        .Y(\PRDATA_0_iv_2_a0[0]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[9]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_807), .C(\PRDATA_0[8] ), .D(N_827), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[13]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_811), .C(\PRDATA_0[8] ), .D(N_831), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[2]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[2]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[2]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[2]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_2_a1[0]  (.A(serdat_0), .B(
        un12_PSELi), .C(un4_PRDATA), .D(CoreAPB3_0_APBmslave0_PSELx), 
        .Y(\PRDATA_0_iv_2_a1[0]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[5]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[5]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[5]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[5]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0[4]  (.A(
        CoreAPB3_0_APBmslave2_PRDATA[4]), .B(
        CoreAPB3_0_APBmslave3_PRDATA[4]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(\PRDATA_0_iv_0[4]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[11]  (.A(PRDATA_regif_sn_N_26), 
        .B(N_809), .C(\PRDATA_0[8] ), .D(N_829), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]));
    
endmodule


module CoreAPB3_Z1(
       iPSELS_0,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR,
       iPSELS_0_0,
       CoreAPB3_0_APBmslave2_PRDATA,
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave0_PRDATA_m_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_1,
       CoreAPB3_0_APBmslave0_PRDATA_m_2,
       CoreAPB3_0_APBmslave1_PRDATA_m,
       CoreAPB3_0_APBmslave4_PRDATA,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       sercon_0,
       sercon_2,
       CoreAPB3_0_APBmslave0_PADDR_0,
       CoreAPB3_0_APBmslave0_PADDR_7,
       serdat_0,
       serdat_2,
       CoreAPB3_0_APBmslave0_PRDATA_m_0_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_4,
       CoreAPB3_0_APBmslave0_PRDATA_m_5,
       CoreAPB3_0_APBmslave0_PRDATA_m_3,
       CoreAPB3_0_APBmslave0_PRDATA_m_2_d0,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_0_APBmslave2_PSELx,
       CoreAPB3_0_APBmslave1_PSELx,
       CoreAPB3_0_APBmslave0_PSELx,
       un4_PRDATA_1,
       controlReg14_3,
       r_N_4_mux,
       un12_PSELi,
       un4_PRDATA,
       un1_PRDATA,
       PRDATA_regif_sn_N_39_mux,
       un14_PRDATA,
       PRDATA_regif_sn_N_26,
       N_809,
       N_829,
       N_810,
       N_830,
       N_807,
       N_827,
       N_808,
       N_828,
       N_812,
       N_832,
       N_806,
       N_826,
       N_813,
       N_833,
       N_811,
       N_831,
       N_840,
       N_842,
       N_837,
       N_841,
       N_839,
       N_838
    );
output [4:4] iPSELS_0;
input  [15:12] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR;
output [4:4] iPSELS_0_0;
input  [7:0] CoreAPB3_0_APBmslave2_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_0;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_1;
input  [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_2;
input  [1:0] CoreAPB3_0_APBmslave1_PRDATA_m;
input  [1:0] CoreAPB3_0_APBmslave4_PRDATA;
output [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
input  sercon_0;
input  sercon_2;
input  CoreAPB3_0_APBmslave0_PADDR_0;
input  CoreAPB3_0_APBmslave0_PADDR_7;
input  serdat_0;
input  serdat_2;
input  CoreAPB3_0_APBmslave0_PRDATA_m_0_d0;
input  CoreAPB3_0_APBmslave0_PRDATA_m_4;
input  CoreAPB3_0_APBmslave0_PRDATA_m_5;
input  CoreAPB3_0_APBmslave0_PRDATA_m_3;
input  CoreAPB3_0_APBmslave0_PRDATA_m_2_d0;
input  mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave3_PSELx;
output CoreAPB3_0_APBmslave2_PSELx;
output CoreAPB3_0_APBmslave1_PSELx;
output CoreAPB3_0_APBmslave0_PSELx;
input  un4_PRDATA_1;
input  controlReg14_3;
output r_N_4_mux;
input  un12_PSELi;
input  un4_PRDATA;
input  un1_PRDATA;
input  PRDATA_regif_sn_N_39_mux;
input  un14_PRDATA;
input  PRDATA_regif_sn_N_26;
input  N_809;
input  N_829;
input  N_810;
input  N_830;
input  N_807;
input  N_827;
input  N_808;
input  N_828;
input  N_812;
input  N_832;
input  N_806;
input  N_826;
input  N_813;
input  N_833;
input  N_811;
input  N_831;
input  N_840;
input  N_842;
input  N_837;
input  N_841;
input  N_839;
input  N_838;

    wire CoreAPB3_0_APBmslave0_PSELx_2, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h1000) )  \iPSELS[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(iPSELS_0[4]), 
        .D(mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave1_PSELx));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h02) )  \iPSELS_0[4]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .C(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .Y(iPSELS_0_0[4])
        );
    CFG4 #( .INIT(16'h0040) )  \iPSELS[2]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(iPSELS_0[4]), 
        .D(mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave2_PSELx));
    COREAPB3_MUXPTOB3 u_mux_p_to_b3 (.CoreAPB3_0_APBmslave2_PRDATA({
        CoreAPB3_0_APBmslave2_PRDATA[7], 
        CoreAPB3_0_APBmslave2_PRDATA[6], 
        CoreAPB3_0_APBmslave2_PRDATA[5], 
        CoreAPB3_0_APBmslave2_PRDATA[4], 
        CoreAPB3_0_APBmslave2_PRDATA[3], 
        CoreAPB3_0_APBmslave2_PRDATA[2], 
        CoreAPB3_0_APBmslave2_PRDATA[1], 
        CoreAPB3_0_APBmslave2_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave3_PRDATA({CoreAPB3_0_APBmslave3_PRDATA[7], 
        CoreAPB3_0_APBmslave3_PRDATA[6], 
        CoreAPB3_0_APBmslave3_PRDATA[5], 
        CoreAPB3_0_APBmslave3_PRDATA[4], 
        CoreAPB3_0_APBmslave3_PRDATA[3], 
        CoreAPB3_0_APBmslave3_PRDATA[2], 
        CoreAPB3_0_APBmslave3_PRDATA[1], 
        CoreAPB3_0_APBmslave3_PRDATA[0]}), .iPSELS_0({iPSELS_0[4]}), 
        .iPSELS_0_0({iPSELS_0_0[4]}), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_0({
        CoreAPB3_0_APBmslave0_PRDATA_m_0[7]}), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_1({
        CoreAPB3_0_APBmslave0_PRDATA_m_1[7]}), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2({
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]}), 
        .CoreAPB3_0_APBmslave1_PRDATA_m({
        CoreAPB3_0_APBmslave1_PRDATA_m[1], 
        CoreAPB3_0_APBmslave1_PRDATA_m[0]}), 
        .CoreAPB3_0_APBmslave4_PRDATA({CoreAPB3_0_APBmslave4_PRDATA[1], 
        CoreAPB3_0_APBmslave4_PRDATA[0]}), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]}), .sercon_0(
        sercon_0), .sercon_2(sercon_2), .CoreAPB3_0_APBmslave0_PADDR_0(
        CoreAPB3_0_APBmslave0_PADDR_0), .CoreAPB3_0_APBmslave0_PADDR_7(
        CoreAPB3_0_APBmslave0_PADDR_7), .serdat_0(serdat_0), .serdat_2(
        serdat_2), .CoreAPB3_0_APBmslave0_PRDATA_m_0_d0(
        CoreAPB3_0_APBmslave0_PRDATA_m_0_d0), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_4(
        CoreAPB3_0_APBmslave0_PRDATA_m_4), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_5(
        CoreAPB3_0_APBmslave0_PRDATA_m_5), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_3(
        CoreAPB3_0_APBmslave0_PRDATA_m_3), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2_d0(
        CoreAPB3_0_APBmslave0_PRDATA_m_2_d0), .un4_PRDATA_1(
        un4_PRDATA_1), .controlReg14_3(controlReg14_3), 
        .CoreAPB3_0_APBmslave0_PSELx(CoreAPB3_0_APBmslave0_PSELx), 
        .r_N_4_mux(r_N_4_mux), .un12_PSELi(un12_PSELi), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_0_APBmslave2_PSELx(CoreAPB3_0_APBmslave2_PSELx), 
        .un4_PRDATA(un4_PRDATA), .un1_PRDATA(un1_PRDATA), 
        .PRDATA_regif_sn_N_39_mux(PRDATA_regif_sn_N_39_mux), 
        .un14_PRDATA(un14_PRDATA), .PRDATA_regif_sn_N_26(
        PRDATA_regif_sn_N_26), .N_809(N_809), .N_829(N_829), .N_810(
        N_810), .N_830(N_830), .N_807(N_807), .N_827(N_827), .N_808(
        N_808), .N_828(N_828), .N_812(N_812), .N_832(N_832), .N_806(
        N_806), .N_826(N_826), .N_813(N_813), .N_833(N_833), .N_811(
        N_811), .N_831(N_831), .N_840(N_840), .N_842(N_842), .N_837(
        N_837), .N_841(N_841), .N_839(N_839), .N_838(N_838));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h1) )  \iPSELS_1[3]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]), .Y(
        CoreAPB3_0_APBmslave0_PSELx_2));
    CFG2 #( .INIT(4'h4) )  \iPSELS_0[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .Y(iPSELS_0[4]));
    CFG4 #( .INIT(16'h8000) )  \iPSELS[3]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .D(
        CoreAPB3_0_APBmslave0_PSELx_2), .Y(CoreAPB3_0_APBmslave3_PSELx)
        );
    CFG4 #( .INIT(16'h0200) )  \iPSELS[0]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .D(
        CoreAPB3_0_APBmslave0_PSELx_2), .Y(CoreAPB3_0_APBmslave0_PSELx)
        );
    
endmodule


module CoreGPIO_Z2(
       GPOUT_reg,
       TRIG_c,
       CoreAPB3_0_APBmslave0_PWDATA,
       ECHO_c,
       CoreAPB3_0_APBmslave0_PADDR,
       gpin3_m_2_0,
       gpin3_m,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       GPOUT_reg40_2,
       GPOUT_reg40,
       un1_WEn_1,
       CoreAPB3_0_APBmslave1_PSELx
    );
output [1:1] GPOUT_reg;
output [0:0] TRIG_c;
input  [1:0] CoreAPB3_0_APBmslave0_PWDATA;
input  [1:1] ECHO_c;
input  [7:0] CoreAPB3_0_APBmslave0_PADDR;
output [1:1] gpin3_m_2_0;
output [1:1] gpin3_m;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output GPOUT_reg40_2;
output GPOUT_reg40;
input  un1_WEn_1;
input  CoreAPB3_0_APBmslave1_PSELx;

    wire VCC_net_1, GPOUT_reg_0_sqmuxa_net_1, GND_net_1, \gpin1[1] , 
        \gpin2[1] , \gpin3[1] , \gpin3_m_1[1] ;
    
    CFG4 #( .INIT(16'h0200) )  
        \xhdl1.GEN_BITS[0].APB_32.GPOUT_reg40_2  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(GPOUT_reg40_2));
    SLE \xhdl1.GEN_BITS[1].gpin1[1]  (.D(ECHO_c[1]), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[1] ));
    CFG4 #( .INIT(16'h8000) )  GPOUT_reg_0_sqmuxa (.A(un1_WEn_1), .B(
        GPOUT_reg40_2), .C(gpin3_m_2_0[1]), .D(
        CoreAPB3_0_APBmslave1_PSELx), .Y(GPOUT_reg_0_sqmuxa_net_1));
    GND GND (.Y(GND_net_1));
    SLE \xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        GPOUT_reg_0_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(GPOUT_reg[1]));
    CFG4 #( .INIT(16'h0001) )  \xhdl1.GEN_BITS[1].gpin3_m_2[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[0]), .D(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(gpin3_m_2_0[1]));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  \xhdl1.GEN_BITS[0].APB_32.GPOUT_reg40  (.A(
        gpin3_m_2_0[1]), .B(GPOUT_reg40_2), .Y(GPOUT_reg40));
    CFG3 #( .INIT(8'h80) )  \xhdl1.GEN_BITS[1].gpin3_RNID0971[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[7]), .B(\gpin3[1] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\gpin3_m_1[1] ));
    SLE \xhdl1.GEN_BITS[1].gpin2[1]  (.D(\gpin1[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin2[1] ));
    SLE \xhdl1.GEN_BITS[1].gpin3[1]  (.D(\gpin2[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin3[1] ));
    CFG4 #( .INIT(16'h1000) )  \xhdl1.GEN_BITS[1].gpin3_RNIBH0T3[1]  (
        .A(CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(\gpin3_m_1[1] ), .D(
        gpin3_m_2_0[1]), .Y(gpin3_m[1]));
    SLE \xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        GPOUT_reg_0_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(TRIG_c[0]));
    
endmodule


module COREI2CREAL_Z4(
       COREI2C_0_0_SDAO_i,
       COREI2C_0_0_SCLO_i,
       COREI2C_0_0_INT,
       CoreAPB3_0_APBmslave0_PADDR,
       CoreAPB3_0_APBmslave0_PRDATA_m_1,
       CoreAPB3_0_APBmslave0_PRDATA_m_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_2,
       TRIG_c,
       gpin3_m_2_0,
       GPOUT_reg,
       gpin3_m,
       CoreAPB3_0_APBmslave1_PRDATA_m,
       CoreAPB3_0_APBmslave0_PWDATA,
       sercon_0,
       sercon_2,
       serdat_2,
       serdat_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_0_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_4,
       CoreAPB3_0_APBmslave0_PRDATA_m_2_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_3,
       CoreAPB3_0_APBmslave0_PRDATA_m_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       r_N_4_mux,
       N_97_1,
       controlReg14_3,
       un4_PRDATA_1,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       un1_WEn_1,
       BIBUF_COREI2C_0_0_SCL_IO_Y,
       BIBUF_COREI2C_0_0_SDA_IO_Y,
       un1_WEn_0,
       un14_PRDATA,
       un1_PRDATA,
       un4_PRDATA,
       CoreAPB3_0_APBmslave0_PSELx,
       un12_PSELi,
       GPOUT_reg40_2,
       CoreAPB3_0_APBmslave1_PSELx,
       GPOUT_reg40
    );
output [0:0] COREI2C_0_0_SDAO_i;
output [0:0] COREI2C_0_0_SCLO_i;
output [0:0] COREI2C_0_0_INT;
input  [8:0] CoreAPB3_0_APBmslave0_PADDR;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_1;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_0;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_2;
input  [0:0] TRIG_c;
input  [1:1] gpin3_m_2_0;
input  [1:1] GPOUT_reg;
input  [1:1] gpin3_m;
output [1:0] CoreAPB3_0_APBmslave1_PRDATA_m;
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output sercon_0;
output sercon_2;
output serdat_2;
output serdat_0;
output CoreAPB3_0_APBmslave0_PRDATA_m_0_d0;
output CoreAPB3_0_APBmslave0_PRDATA_m_4;
output CoreAPB3_0_APBmslave0_PRDATA_m_2_d0;
output CoreAPB3_0_APBmslave0_PRDATA_m_3;
output CoreAPB3_0_APBmslave0_PRDATA_m_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  r_N_4_mux;
output N_97_1;
output controlReg14_3;
output un4_PRDATA_1;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
output un1_WEn_1;
input  BIBUF_COREI2C_0_0_SCL_IO_Y;
input  BIBUF_COREI2C_0_0_SDA_IO_Y;
output un1_WEn_0;
output un14_PRDATA;
output un1_PRDATA;
output un4_PRDATA;
input  CoreAPB3_0_APBmslave0_PSELx;
input  un12_PSELi;
input  GPOUT_reg40_2;
input  CoreAPB3_0_APBmslave1_PSELx;
input  GPOUT_reg40;

    wire \COREI2C_0_0_SDAO[0] , \COREI2C_0_0_SCLO[0] , 
        \fsmdet[3]_net_1 , \fsmdet_i_0[3] , SCLInt_net_1, SCLInt_i_0, 
        \SDAI_ff_reg[3]_net_1 , GND_net_1, N_68_i_0, VCC_net_1, 
        \SCLI_ff_reg[0]_net_1 , \SCLI_ff_reg_3[0] , 
        \SCLI_ff_reg[1]_net_1 , N_293_i_0, \SCLI_ff_reg[2]_net_1 , 
        N_294_i_0, \SCLI_ff_reg[3]_net_1 , N_295_i_0, 
        \SDAI_ff_reg[0]_net_1 , \SDAI_ff_reg_3[0] , 
        \SDAI_ff_reg[1]_net_1 , N_64_i_0, \SDAI_ff_reg[2]_net_1 , 
        N_66_i_0, \sercon[7]_net_1 , sercon18, \PCLK_count2[0]_net_1 , 
        \PCLK_count2_4[0]_net_1 , \PCLK_count2[1]_net_1 , 
        \PCLK_count2_4[1]_net_1 , \framesync[0]_net_1 , 
        \framesync_6[0] , \framesync[1]_net_1 , \framesync_6[1] , 
        \framesync[2]_net_1 , \framesync_6[2] , \framesync[3]_net_1 , 
        \framesync_6[3] , \PCLK_count1[0]_net_1 , N_340_i_0, 
        \PCLK_count1[1]_net_1 , N_341_i_0, \PCLK_count1[2]_net_1 , 
        N_342_i_0, \PCLK_count1[3]_net_1 , \PCLK_count1_4[3] , 
        \indelay[0]_net_1 , \indelay_4[0]_net_1 , \indelay[1]_net_1 , 
        \indelay_4[1]_net_1 , \indelay[2]_net_1 , \indelay_4[2]_net_1 , 
        \sercon[1]_net_1 , \sercon_9[3] , \sercon[4]_net_1 , N_62_i_0, 
        \sercon[5]_net_1 , \sercon[6]_net_1 , \serdat[1]_net_1 , 
        \serdat_19[1] , un1_N_9_mux_i_0, \serdat_19[2] , 
        \serdat[3]_net_1 , \serdat_19[3] , \serdat[4]_net_1 , 
        \serdat_19[4] , \serdat[5]_net_1 , \serdat_19[5] , 
        \serdat[6]_net_1 , \serdat_19[6] , \serdat[7]_net_1 , 
        \serdat_19[7] , \serdat_19[0] , \sersta[4]_net_1 , 
        \sersta_3[4] , sclscl_net_1, \fsmmod[5]_net_1 , 
        sclscl_1_sqmuxa_i_0, SDAInt_net_1, un1_SDAInt5, un1_SCLInt5, 
        nedetect_net_1, nedetect_0_sqmuxa, pedetect_0_sqmuxa_3, 
        starto_en_net_1, N_344, starto_en_1_sqmuxa_i_0_net_1, 
        pedetect_net_1, pedetect_0_sqmuxa, N_262, \fsmsta[0]_net_1 , 
        \fsmsta_9[0] , un1_ens1_pre_1_sqmuxa_i_0_net_1, 
        \fsmsta[1]_net_1 , N_1328_i_0, \fsmsta[2]_net_1 , 
        \fsmsta_9[2] , \fsmsta[3]_net_1 , N_94, \fsmsta[4]_net_1 , 
        \fsmsta_9[4] , \sersta[0]_net_1 , \sersta_3[0] , 
        \sersta[1]_net_1 , \sersta_3[1] , \sersta[2]_net_1 , 
        \sersta_3[2] , \sersta[3]_net_1 , \sersta_3[3] , ack_net_1, 
        ack_10, N_1272, SDAO_int_1_sqmuxa_i_0, bsd7_net_1, 
        bsd7_10_iv_i_0, bsd7_tmp_net_1, bsd7_tmp_7, adrcomp_net_1, 
        un1_adrcomp14_1, adrcomp_2_sqmuxa_i_0, ack_bit_net_1, 
        ack_bit_1_sqmuxa_net_1, PCLKint_net_1, PCLKint_4, 
        un1_fsmdet_1_i_0, busfree_net_1, un1_fsmdet, adrcompen_net_1, 
        un1_adrcomp14_net_1, adrcompen_2_sqmuxa_i_0, \fsmdet[0]_net_1 , 
        \fsmdet[1]_net_1 , N_871_i_0, \fsmdet[2]_net_1 , N_873_i_0, 
        N_875_i_0, \fsmdet[4]_net_1 , N_877_i_0, \fsmdet[5]_net_1 , 
        N_879_i_0, \fsmdet[6]_net_1 , N_881_i_0, \fsmsync[0]_net_1 , 
        \fsmsync_ns[0] , \fsmsync[1]_net_1 , N_955_i_0, 
        \fsmsync[2]_net_1 , N_957_i_0, \fsmsync[3]_net_1 , N_959_i_0, 
        \fsmsync[4]_net_1 , N_961_i_0, \fsmsync[5]_net_1 , N_963_i_0, 
        \fsmsync[6]_net_1 , N_965_i_0, \fsmmod[0]_net_1 , 
        \fsmmod_ns[0] , \fsmmod[1]_net_1 , \fsmmod_ns[1] , 
        \fsmmod[2]_net_1 , N_1010_i_0, \fsmmod[3]_net_1 , 
        \fsmmod_ns[3] , \fsmmod[4]_net_1 , N_1013_i_0, \fsmmod_ns[5] , 
        \fsmmod[6]_net_1 , N_1016_i_0, PCLK_count1_ov_net_1, 
        PCLK_count1_ov_3, PCLKint_ff_net_1, PCLKint_ff_3, 
        PCLK_count2_ov_net_1, PCLK_count2_ov_0_sqmuxa_net_1, 
        SCLO_int5_i_0, un1_framesync_2, CO1, counter_PRESETN_net_1, 
        CO0, N_220, N_980, N_129, counter_PRESETN_1, 
        counter_PRESETN_0_net_1, N_490, \fsmsta_9_0_o2_1_2_1[0] , 
        N_400, \fsmsta_9_0_o2_1_1[0] , N_353, N_412, N_543, N_359, 
        N_404, fsmsta_9_0_372_i_0_a2_3_1, N_444, 
        fsmsta_9_0_372_i_0_o2_6_0, N_480, framesync24, N_554, 
        \fsmsta_9_0_a2_4_0[0] , N_443, N_527, 
        un1_ens1_pre_1_sqmuxa_i_0_1_net_1, N_514, N_380, 
        \fsmsta_9_0_1_1[0] , \fsmsta_9_0_1[0] , un1_framesync24, N_370, 
        N_355, \fsmmod_ns_0_0_o2_1[3]_net_1 , N_162, adrcomp12, 
        adrcomp7_0_0, adrcomp_2_sqmuxa_0_1_net_1, sersta77_2, N_360, 
        N_358, fsmsta_9_0_372_i_0_a2_0_1, fsmsta_9_0_372_i_0_a2_0_0, 
        N_356, N_441, \fsmsta_9_0_o2_6_1_1[0] , \fsmsta_9_0_o2_6_1[0] , 
        N_365, \fsmsta_9_0_m2_bm[2] , \fsmsta_9_0_m2_am[2] , N_226, 
        bsd7_tmp_7_sm0, bsd7_tmp_7_am, bsd7_tmp_7_bm, un1_sersta65_1_0, 
        N_1236, un1_sersta65_1_1, un1_sersta65_1, d_N_5_mux, 
        bsd7_N_12_mux, bsd7_i_m, un1_sercon_1_6, un1_sersta64_1, N_548, 
        N_479, N_394, \fsmmod_ns_0_0_a2_0[5]_net_1 , 
        \fsmmod_ns_0_0_a2_0_0[5]_net_1 , \fsmsta_9_0_a2_2_0[4] , 
        \fsmsync_ns_0_a3_0_1[0]_net_1 , \fsmsta_9_0_o2_3_0[2] , 
        un12_PSELi_0, N_492, N_531, N_438_1, N_155, fsmsync_nxt35, 
        N_361, N_140_i, N_393, N_372, bsd7_tmp_i_m_1, N_1028_2, N_526, 
        N_364, N_367, N_416, PRDATA_N_9, r_N_3_0, SDAO_int_6_0_312_1, 
        bsd7_10_iv_1_a0_2, SDAO_int_1_sqmuxa_1_net_1, 
        \PCLK_count1_4_0_a2_0_0[3] , un1_fsmsync_2, bsd7_m6_0, 
        sercon_m2_e_2_1, sercon_m2_e_3_1, sercon_m2_e_0_1, 
        sercon_m2_e_1, un14_PRDATA_0_net_1, un9_PRDATA_1_net_1, 
        un1_sercon_1_3, \fsmsta_9_0_a2_3_1[4] , 
        fsmsta_9_2_342_i_i_a2_10_0, \fsmmod_ns_i_0_a2_0_0[2]_net_1 , 
        fsmsta_9_0_372_i_0_a2_12_0, \fsmsta_9_0_a2_8_0[2] , N_510, 
        N_512, N_827, un18_counter_PRESETN_net_1, un1_ack_1_0, N_244, 
        framesync_6_e2_1, un1_framesync_1, un14_counter_PRESETN_net_1, 
        fsmsta_m2_e_0, N_1235, N_549, N_979, N_407, N_507, N_504, 
        N_289, N_524, N_374, N_547, N_185, SDAO_int6, N_533, N_401, 
        N_224, N_221, SDAO_int_6_0_312_a5_0, bsd7_10_iv_1_a0_3, 
        un1_PSEL_0, \fsmmod_ns_0_0_a2_1[3] , SDAO_int_1_sqmuxa_3_net_1, 
        fsmsta_9_2_342_i_i_o2_3_0, un1_sercon_1_5, \sersta_3_0_1[3] , 
        fsmsta_9_2_342_i_i_a2_8_0, fsmsta_9_0_372_i_0_o2_11_0, 
        un1_fsmdet_1_2_net_1, \fsmmod_ns_i_0_a2_0_2[2]_net_1 , 
        \fsmsta_9_0_a2_2_2[4] , \fsmsta_9_0_a2_0_1[4] , 
        un1_framesync24_1, \sercon_m[4] , \sercon_m[3] , N_496, N_985, 
        N_471, N_474, N_499, N_200, N_476, N_460, N_418, \sercon_m[6] , 
        \sercon_m[1] , \serdat_m[1] , N_994, N_466, N_385, N_497, 
        N_438, N_292, N_291, N_477, un1_sersta58, N_213, un1_nedetect, 
        N_452, N_542, \serdat_RNI49U42[5]_net_1 , N_414, N_410, 
        un1_sersta58_0, N_384, SDAO_int_1_sqmuxa_4_net_1, 
        \fsmmod_ns_i_0_0[4]_net_1 , \fsmmod_ns_0_0_0[0]_net_1 , 
        bsd7_m6_3, fsmsta_9_0_372_i_0_o2_1_1, 
        \fsmsync_ns_i_0[6]_net_1 , \fsmsta_9_0_o2_1_2[2] , 
        \fsmsta_9_0_o2_1_0[2] , \fsmsync_ns_i_0[2]_net_1 , 
        \fsmsync_ns_i_0[3]_net_1 , \fsmsta_9_0_a2_1_2[4] , 
        \sersta_3_0_1[1] , fsmsta_9_0_372_i_0_o2_12_1, 
        \sercon_9_0_a2_0_1[3] , N_990, N_972, N_255, framesync14, 
        framesync10, N_455, N_453, N_152, N_151, N_973, N_509, N_317, 
        N_395, N_480_2, bsd7_tmp_i_m_1_0, \serdat_i_m_3_1[7] , 
        \PRDATA_0_iv_0[4]_net_1 , \PRDATA_0_iv_0[3]_net_1 , 
        \PRDATA_0_iv_0[6]_net_1 , \fsmsta_9_0_0[4] , 
        \sercon_9_0_0_a1_tz_0[3] , fsmsta_9_0_372_i_0_o2_1_3, 
        \fsmsync_ns_i_1[6]_net_1 , \fsmsta_9_0_o2_1_3[2] , 
        \fsmsync_ns_0_1[0]_net_1 , bsd7_10_iv_1_a0_2_RNI6O401, 
        un1_sersta69, N_555, N_301, N_1288, \sercon_9_0_0_a0[3] , 
        N_530, serdat4, N_227, N_419, N_447, \PWDATA_i_m_1[7] , 
        \fsmsta_9_0_o2_3_0[0] , serdat_2_sqmuxa_out, 
        \fsmmod_ns_0_0_0[5]_net_1 , \fsmsta_9_0_1[4] , 
        fsmsta_9_2_342_i_i_o2_3_2, fsmsta_9_0_372_i_0_o2_1_4, 
        \fsmsta_9_0_o2_1_4[2] , N_551, N_238, N_398, N_228, 
        framesync_6_e2, CO2, \serdat_i_m_3_0_0[7] , m3_0, 
        bsd7_10_iv_1_a1, ack_10_u_yy, ack_10_u_xx, 
        fsmsta_9_2_342_i_i_0, fsmsta_9_0_372_i_0_2, 
        fsmsta_9_2_342_i_i_o2_0, N_298, \framesync_6_m2[3] , 
        un1_sersta65, serdat48, bsd7_10_iv_1, fsmsta_9_0_372_i_0_4, 
        fsmsta_9_0_372_i_0_3, \fsmsta_9_0_3[4] , N_413, N_297, 
        N_2_4_tz, ack_1_sqmuxa_1_net_1, N_442, N_1289, 
        \fsmsta_9_RNO[0] , N_449, serdat_1_sqmuxa_1_net_1, 
        un1_serdat_2_sqmuxa_1_tz, \sercon_9_0_0[3] , N_117;
    
    CFG4 #( .INIT(16'hF080) )  \PRDATA_0_iv_0_RNISGIF1[3]  (.A(
        un4_PRDATA), .B(\serdat[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]), .D(
        \PRDATA_0_iv_0[3]_net_1 ), .Y(
        CoreAPB3_0_APBmslave0_PRDATA_m_2_d0));
    CFG4 #( .INIT(16'hF3A3) )  \fsmsta_sync_proc.fsmsta_9_0_m2[4]  (.A(
        \fsmmod[6]_net_1 ), .B(\fsmdet[5]_net_1 ), .C(
        \fsmdet[3]_net_1 ), .D(\fsmmod[1]_net_1 ), .Y(N_221));
    CFG3 #( .INIT(8'h54) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_12_0  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[4]_net_1 ), .Y(fsmsta_9_0_372_i_0_a2_12_0));
    CFG2 #( .INIT(4'hB) )  \PCLKint_write_proc.PCLKint_4  (.A(
        counter_PRESETN_net_1), .B(PCLKint_net_1), .Y(PCLKint_4));
    CFG4 #( .INIT(16'h0105) )  \serdat_write_proc.bsd7_10_iv_i  (.A(
        bsd7_10_iv_1), .B(\PWDATA_i_m_1[7] ), .C(bsd7_i_m), .D(serdat4)
        , .Y(bsd7_10_iv_i_0));
    SLE \sercon[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[1]_net_1 ));
    CFG4 #( .INIT(16'hFFD0) )  ack_RNO_0 (.A(un1_sersta65), .B(
        ack_1_sqmuxa_1_net_1), .C(pedetect_net_1), .D(
        serdat_2_sqmuxa_out), .Y(un1_serdat_2_sqmuxa_1_tz));
    CFG4 #( .INIT(16'h8000) )  \sercon_write_proc.sercon18  (.A(
        un12_PSELi), .B(un1_WEn_1), .C(CoreAPB3_0_APBmslave0_PSELx), 
        .D(un1_PRDATA), .Y(sercon18));
    CFG4 #( .INIT(16'h0F0E) )  \fsmsta_sync_proc.fsmsta_9_RNO[0]  (.A(
        N_400), .B(N_412), .C(counter_PRESETN_1), .D(N_543), .Y(
        \fsmsta_9_RNO[0] ));
    CFG4 #( .INIT(16'h5554) )  \sercon_write_proc.un1_framesync24_1  (
        .A(\framesync[3]_net_1 ), .B(\framesync[0]_net_1 ), .C(
        \framesync[2]_net_1 ), .D(\framesync[1]_net_1 ), .Y(
        un1_framesync24_1));
    CFG4 #( .INIT(16'h0008) )  \sercon_write_proc.un1_PSEL_0_0  (.A(
        un1_WEn_1), .B(un12_PSELi_0), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(un1_PSEL_0));
    CFG2 #( .INIT(4'h8) )  \un1_framesync_1_1.CO2  (.A(CO1), .B(
        \framesync[2]_net_1 ), .Y(CO2));
    CFG4 #( .INIT(16'hFFFE) )  un1_ens1_pre_1_sqmuxa_i_0 (.A(N_443), 
        .B(N_527), .C(un1_ens1_pre_1_sqmuxa_i_0_1_net_1), .D(N_514), 
        .Y(un1_ens1_pre_1_sqmuxa_i_0_net_1));
    CFG4 #( .INIT(16'h01A1) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_9  (.A(
        \fsmsta[4]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(N_358), .D(
        \fsmsta_9_0_o2_3_0[2] ), .Y(N_151));
    CFG4 #( .INIT(16'hEEE2) )  \fsmsta_sync_proc.fsmsta_9_0_m2_bm[2]  
        (.A(N_555), .B(N_129), .C(\fsmsta_9_0_o2_1_3[2] ), .D(
        \fsmsta_9_0_o2_1_4[2] ), .Y(\fsmsta_9_0_m2_bm[2] ));
    CFG4 #( .INIT(16'h2202) )  \fsmsta_sync_proc.fsmsta_9_0_a2_17[0]  
        (.A(SDAInt_net_1), .B(\fsmsta[3]_net_1 ), .C(\fsmsta[1]_net_1 )
        , .D(\fsmsta[4]_net_1 ), .Y(N_510));
    SLE \fsmdet[1]  (.D(N_871_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[1]_net_1 ));
    CFG4 #( .INIT(16'h3ACA) )  
        \framesync_write_proc.framesync_6_enl[2]  (.A(
        \fsmdet[3]_net_1 ), .B(\framesync[2]_net_1 ), .C(
        framesync_6_e2), .D(CO1), .Y(\framesync_6[2] ));
    SLE SDAInt (.D(\SDAI_ff_reg[0]_net_1 ), .CLK(GL0_INST), .EN(
        un1_SDAInt5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        SDAInt_net_1));
    SLE starto_en (.D(N_344), .CLK(GL0_INST), .EN(
        starto_en_1_sqmuxa_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(starto_en_net_1));
    CFG1 #( .INIT(2'h1) )  SDAO_int_RNINGI9 (.A(\COREI2C_0_0_SDAO[0] ), 
        .Y(COREI2C_0_0_SDAO_i[0]));
    CFG4 #( .INIT(16'h8000) )  
        \serdat_write_proc.bsd7_10_iv_1_a0_2_RNI6O401  (.A(
        bsd7_10_iv_1_a0_2), .B(un12_PSELi_0), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(un4_PRDATA), .Y(
        bsd7_10_iv_1_a0_2_RNI6O401));
    SLE \serdat[4]  (.D(\serdat_19[4] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[4]_net_1 ));
    CFG4 #( .INIT(16'h1110) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_a2_0  (.A(adrcomp_net_1), 
        .B(\fsmdet[3]_net_1 ), .C(N_395), .D(N_413), .Y(N_449));
    SLE \fsmsta[4]  (.D(\fsmsta_9[4] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fsmsta[4]_net_1 ));
    SLE \SCLI_ff_reg[1]  (.D(N_293_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[1]_net_1 ));
    SLE pedetect (.D(pedetect_0_sqmuxa), .CLK(GL0_INST), .EN(N_262), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(pedetect_net_1)
        );
    CFG2 #( .INIT(4'hD) )  \fsmmod_ns_i_0_o2_0[6]  (.A(
        \sercon[6]_net_1 ), .B(\fsmdet[5]_net_1 ), .Y(N_372));
    SLE \fsmmod[4]  (.D(N_1013_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[4]_net_1 ));
    CFG4 #( .INIT(16'hFFFB) )  \busfree_write_proc.un1_fsmdet_0  (.A(
        counter_PRESETN_1), .B(\sercon[6]_net_1 ), .C(N_548), .D(
        adrcomp12), .Y(un1_fsmdet));
    CFG4 #( .INIT(16'hFFF2) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_1_4  (.A(N_533), .B(
        \COREI2C_0_0_SDAO[0] ), .C(fsmsta_9_0_372_i_0_o2_1_3), .D(
        N_499), .Y(fsmsta_9_0_372_i_0_o2_1_4));
    CFG2 #( .INIT(4'h1) )  \fsmsync_ns_0_a3_0_1[0]  (.A(
        \fsmmod[4]_net_1 ), .B(\fsmmod[3]_net_1 ), .Y(
        \fsmsync_ns_0_a3_0_1[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \fsmmod_ns_0_0_a2_1[0]  (.A(N_547), .B(
        \fsmmod[4]_net_1 ), .Y(N_548));
    CFG4 #( .INIT(16'hFFF8) )  \fsmmod_ns_0_0[0]  (.A(
        \fsmmod[0]_net_1 ), .B(N_200), .C(\fsmmod_ns_0_0_0[0]_net_1 ), 
        .D(N_398), .Y(\fsmmod_ns[0] ));
    CFG2 #( .INIT(4'hE) )  counter_PRESETN_1_0_o2 (.A(
        \fsmdet[3]_net_1 ), .B(\fsmdet[5]_net_1 ), .Y(
        counter_PRESETN_1));
    SLE ack (.D(ack_10), .CLK(GL0_INST), .EN(\sercon[6]_net_1 ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(ack_net_1));
    CFG4 #( .INIT(16'h0004) )  \serdat_write_proc.bsd7_10_iv_i_RNO_3  
        (.A(CoreAPB3_0_APBmslave0_PADDR[8]), .B(bsd7_m6_0), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(bsd7_m6_3));
    CFG4 #( .INIT(16'hEFEE) )  \fsmsta_sync_proc.fsmsta_9_0_o2_6[0]  (
        .A(\fsmsta_9_0_o2_6_1[0] ), .B(N_530), .C(N_356), .D(N_385), 
        .Y(N_412));
    SLE \fsmsta[3]  (.D(N_94), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fsmsta[3]_net_1 ));
    CFG4 #( .INIT(16'h020E) )  \PCLK_counter1_proc.PCLK_count1_4_0[3]  
        (.A(\PCLK_count1_4_0_a2_0_0[3] ), .B(\PCLK_count1[3]_net_1 ), 
        .C(counter_PRESETN_net_1), .D(N_220), .Y(\PCLK_count1_4[3] ));
    CFG3 #( .INIT(8'h01) )  \framesync_write_proc.framesync_6_e2_1  (
        .A(\fsmdet[5]_net_1 ), .B(\fsmdet[3]_net_1 ), .C(
        bsd7_tmp_i_m_1), .Y(framesync_6_e2_1));
    SLE \serdat[2]  (.D(\serdat_19[2] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(serdat_2));
    CFG3 #( .INIT(8'h01) )  un9_PRDATA_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[1]), .C(
        CoreAPB3_0_APBmslave0_PADDR[0]), .Y(un9_PRDATA_1_net_1));
    CFG4 #( .INIT(16'hF080) )  \PRDATA_0_iv_0_RNIUIIF1[4]  (.A(
        un4_PRDATA), .B(\serdat[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]), .D(
        \PRDATA_0_iv_0[4]_net_1 ), .Y(CoreAPB3_0_APBmslave0_PRDATA_m_3)
        );
    CFG4 #( .INIT(16'h5556) )  \sercon_write_proc.un1_framesync24  (.A(
        \framesync[3]_net_1 ), .B(\framesync[0]_net_1 ), .C(
        \framesync[2]_net_1 ), .D(\framesync[1]_net_1 ), .Y(
        un1_framesync24));
    CFG3 #( .INIT(8'hF4) )  \fsmsta_sync_proc.fsmsta_9_0_o2_12[0]  (.A(
        \COREI2C_0_0_SDAO[0] ), .B(N_492), .C(N_510), .Y(N_385));
    CFG3 #( .INIT(8'h08) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_15  (.A(
        \fsmsta[3]_net_1 ), .B(N_480_2), .C(\COREI2C_0_0_SDAO[0] ), .Y(
        N_480));
    CFG3 #( .INIT(8'h08) )  \serdat_write_proc.bsd7_10_iv_1_a1_RNO  (
        .A(bsd7_tmp_i_m_1), .B(un1_sersta58_0), .C(bsd7_tmp_net_1), .Y(
        bsd7_tmp_i_m_1_0));
    CFG3 #( .INIT(8'hF2) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1_1[2]  (
        .A(\fsmsta_9_0_a2_8_0[2] ), .B(N_355), .C(N_474), .Y(
        \fsmsta_9_0_o2_1_0[2] ));
    CFG3 #( .INIT(8'h20) )  starto_en_1_sqmuxa_i_0_1 (.A(SCLInt_net_1), 
        .B(\fsmmod[5]_net_1 ), .C(busfree_net_1), .Y(N_344));
    CFG4 #( .INIT(16'hFFFD) )  \fsmsync_ns_0_o3_0[0]  (.A(
        PCLKint_net_1), .B(N_438), .C(\fsmmod[4]_net_1 ), .D(
        PCLKint_ff_net_1), .Y(N_972));
    CFG4 #( .INIT(16'h1000) )  \fsmsync_ns_0_a3_0[0]  (.A(
        \fsmmod[1]_net_1 ), .B(\fsmmod[2]_net_1 ), .C(N_438_1), .D(
        \fsmsync_ns_0_a3_0_1[0]_net_1 ), .Y(N_985));
    CFG4 #( .INIT(16'hA020) )  \fsmsta_sync_proc.fsmsta_9_0_a2_4[2]  (
        .A(sersta77_2), .B(N_358), .C(\fsmsta[2]_net_1 ), .D(
        \fsmsta_9_0_o2_3_0[2] ), .Y(N_471));
    CFG3 #( .INIT(8'h31) )  \fsmmod_ns_i_0_a2[6]  (.A(
        \fsmmod[3]_net_1 ), .B(\fsmmod[6]_net_1 ), .C(N_407), .Y(N_317)
        );
    CFG2 #( .INIT(4'h7) )  \sersta_write_proc.sersta_3_0_o2[3]  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_416));
    CFG4 #( .INIT(16'h1230) )  \PCLK_count1_RNO[2]  (.A(
        \PCLK_count1[0]_net_1 ), .B(N_238), .C(\PCLK_count1[2]_net_1 ), 
        .D(\PCLK_count1[1]_net_1 ), .Y(N_342_i_0));
    CFG2 #( .INIT(4'hE) )  \framesync_write_proc.un1_nedetect  (.A(
        un1_framesync_2), .B(nedetect_net_1), .Y(un1_nedetect));
    CFG4 #( .INIT(16'h0020) )  SDAO_int_1_sqmuxa_4 (.A(
        \sercon[6]_net_1 ), .B(\fsmmod[3]_net_1 ), .C(
        SDAO_int_1_sqmuxa_3_net_1), .D(SDAO_int6), .Y(
        SDAO_int_1_sqmuxa_4_net_1));
    CFG4 #( .INIT(16'hECCC) )  \PRDATA_0_iv_0[6]  (.A(N_97_1), .B(
        \sercon_m[6] ), .C(\sersta[3]_net_1 ), .D(un9_PRDATA_1_net_1), 
        .Y(\PRDATA_0_iv_0[6]_net_1 ));
    CFG4 #( .INIT(16'h4EE4) )  
        \framesync_write_proc.framesync_6_enl[3]  (.A(framesync_6_e2), 
        .B(\framesync_6_m2[3] ), .C(\framesync[3]_net_1 ), .D(CO2), .Y(
        \framesync_6[3] ));
    CFG4 #( .INIT(16'h0CAE) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1_3[2]  
        (.A(N_524), .B(N_1236), .C(\COREI2C_0_0_SDAO[0] ), .D(
        \fsmsta[1]_net_1 ), .Y(\fsmsta_9_0_o2_1_2[2] ));
    CFG2 #( .INIT(4'hE) )  \PCLK_counter1_proc.PCLK_count1_4_i_o2[0]  
        (.A(\PCLK_count1[1]_net_1 ), .B(\PCLK_count1[2]_net_1 ), .Y(
        N_155));
    CFG2 #( .INIT(4'h1) )  \serdat_write_proc.un4_PRDATA_2_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(controlReg14_3));
    CFG4 #( .INIT(16'h4044) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_3  (.A(
        counter_PRESETN_1), .B(N_359), .C(N_404), .D(
        fsmsta_9_0_372_i_0_a2_3_1), .Y(N_444));
    CFG3 #( .INIT(8'h10) )  un14_PRDATA_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(un14_PRDATA_0_net_1), .Y(
        un14_PRDATA));
    CFG4 #( .INIT(16'h1000) )  \SDAO_int_write_proc.un1_framesync_2  (
        .A(\framesync[2]_net_1 ), .B(\framesync[1]_net_1 ), .C(
        \framesync[0]_net_1 ), .D(\framesync[3]_net_1 ), .Y(
        un1_framesync_2));
    CFG2 #( .INIT(4'h1) )  pedetect_0_sqmuxa_0_a2 (.A(
        pedetect_0_sqmuxa_3), .B(SCLInt_net_1), .Y(pedetect_0_sqmuxa));
    CFG4 #( .INIT(16'hCCDC) )  \fsmmod_ns_0_0[5]  (.A(N_398), .B(
        \fsmmod_ns_0_0_0[5]_net_1 ), .C(\fsmmod_ns_0_0_a2_0[5]_net_1 ), 
        .D(N_200), .Y(\fsmmod_ns[5] ));
    SLE \fsmmod[3]  (.D(\fsmmod_ns[3] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \framesync_write_proc.framesync14_0_a2  (.A(
        N_533), .B(\fsmsta[0]_net_1 ), .Y(N_466));
    CFG4 #( .INIT(16'hAEFF) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_o4_0  (.A(bsd7_net_1), 
        .B(\framesync[3]_net_1 ), .C(un1_framesync_2), .D(
        un1_sersta58_0), .Y(N_1288));
    CFG4 #( .INIT(16'h0200) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_6  (.A(ack_net_1), .B(
        \fsmsta[2]_net_1 ), .C(counter_PRESETN_1), .D(N_542), .Y(N_447)
        );
    CFG4 #( .INIT(16'h1050) )  \framesync_write_proc.framesync_6_e2  (
        .A(un1_framesync_2), .B(nedetect_net_1), .C(framesync_6_e2_1), 
        .D(framesync24), .Y(framesync_6_e2));
    CFG4 #( .INIT(16'h8000) )  \adrcomp_write_proc.un1_sercon_1_3  (.A(
        \serdat[6]_net_1 ), .B(sercon_2), .C(adrcompen_net_1), .D(
        \serdat[1]_net_1 ), .Y(un1_sercon_1_3));
    CFG3 #( .INIT(8'h54) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_11_0  (.A(
        \fsmsta[1]_net_1 ), .B(N_367), .C(\fsmsta[3]_net_1 ), .Y(
        fsmsta_9_0_372_i_0_o2_11_0));
    CFG4 #( .INIT(16'h2000) )  \adrcomp_write_proc.un1_sercon_1_6  (.A(
        nedetect_net_1), .B(\serdat[5]_net_1 ), .C(un1_sercon_1_5), .D(
        un1_sercon_1_3), .Y(un1_sercon_1_6));
    CFG4 #( .INIT(16'hFFFE) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_2  
        (.A(N_443), .B(N_527), .C(N_441), .D(N_447), .Y(
        fsmsta_9_0_372_i_0_2));
    CFG3 #( .INIT(8'hAE) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_12  (.A(
        fsmsta_9_0_372_i_0_o2_12_1), .B(\fsmsta[2]_net_1 ), .C(N_360), 
        .Y(N_555));
    CFG3 #( .INIT(8'hAE) )  \serdat_write_proc.bsd7_tmp_7_am_RNO  (.A(
        bsd7_tmp_net_1), .B(\serdat_i_m_3_1[7] ), .C(un4_PRDATA), .Y(
        \serdat_i_m_3_0_0[7] ));
    SLE \serdat[7]  (.D(\serdat_19[7] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[7]_net_1 ));
    SLE \sercon[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(sercon_2));
    CFG3 #( .INIT(8'hC4) )  \fsmsta_sync_proc.fsmsta_9_0_a2_0[2]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(N_361), .Y(N_477)
        );
    CFG4 #( .INIT(16'hFFFE) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_11  (.A(N_533), .B(
        N_524), .C(fsmsta_9_0_372_i_0_o2_11_0), .D(N_527), .Y(N_554));
    CFG4 #( .INIT(16'hFFCA) )  \fsmsta_sync_proc.fsmsta_9[0]  (.A(
        \fsmsta_9_RNO[0] ), .B(N_353), .C(fsmsta_m2_e_0), .D(
        \fsmsta_9_0_1[0] ), .Y(\fsmsta_9[0] ));
    CFG4 #( .INIT(16'h1555) )  \serdat_write_proc.bsd7_10_iv_0  (.A(
        bsd7_10_iv_1_a1), .B(un4_PRDATA), .C(bsd7_10_iv_1_a0_3), .D(
        CoreAPB3_0_APBmslave0_PSELx), .Y(bsd7_10_iv_1));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h02) )  \serdat_write_proc.serdat48  (.A(
        un1_sersta65_1), .B(\fsmdet[3]_net_1 ), .C(un1_sersta58_0), .Y(
        serdat48));
    CFG4 #( .INIT(16'hFFFE) )  counter_PRESETN_0 (.A(
        \fsmsync[1]_net_1 ), .B(\fsmsync[4]_net_1 ), .C(
        \fsmsync[5]_net_1 ), .D(counter_PRESETN_1), .Y(
        counter_PRESETN_0_net_1));
    SLE sclscl (.D(\fsmmod[5]_net_1 ), .CLK(GL0_INST), .EN(
        sclscl_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sclscl_net_1));
    CFG2 #( .INIT(4'h8) )  \sersta_write_proc.sersta_3_0_a2_0[4]  (.A(
        N_549), .B(\fsmsta[3]_net_1 ), .Y(N_292));
    CFG4 #( .INIT(16'hEEE4) )  PRDATA_m6_0_m4_RNIL47A1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(PRDATA_N_9), .C(
        \serdat[7]_net_1 ), .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        CoreAPB3_0_APBmslave0_PRDATA_m_0[7]));
    CFG3 #( .INIT(8'h12) )  \PCLK_count2_4[0]  (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN_net_1), .C(
        \PCLK_count2[0]_net_1 ), .Y(\PCLK_count2_4[0]_net_1 ));
    CFG4 #( .INIT(16'h055D) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_0_1  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \COREI2C_0_0_SDAO[0] ), .D(\fsmsta[0]_net_1 ), .Y(
        fsmsta_9_0_372_i_0_a2_0_1));
    CFG3 #( .INIT(8'h04) )  \framesync_write_proc.framesync10  (.A(
        COREI2C_0_0_INT[0]), .B(un1_sersta58), .C(\sercon[4]_net_1 ), 
        .Y(framesync10));
    CFG1 #( .INIT(2'h1) )  busfree_RNO (.A(\fsmdet[3]_net_1 ), .Y(
        \fsmdet_i_0[3] ));
    SLE \SCLI_ff_reg[0]  (.D(\SCLI_ff_reg_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[0]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2  (
        .A(adrcomp_net_1), .B(adrcompen_net_1), .Y(N_359));
    CFG4 #( .INIT(16'hFFDF) )  \fsmsta_sync_proc.fsmsta_9_0_o2_3[4]  (
        .A(\fsmsta[2]_net_1 ), .B(N_1028_2), .C(\framesync[3]_net_1 ), 
        .D(\framesync[0]_net_1 ), .Y(N_356));
    CFG4 #( .INIT(16'h202F) )  \serdat_RNI49U42[5]  (.A(
        \serdat[5]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .D(r_N_3_0), .Y(
        \serdat_RNI49U42[5]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \fsmsync_RNO[6]  (.A(\fsmsync[6]_net_1 )
        , .B(\sercon[4]_net_1 ), .C(N_973), .D(
        \fsmsync_ns_i_1[6]_net_1 ), .Y(N_965_i_0));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_proc.SDAI_ff_reg_3[0]  (.A(
        \sercon[6]_net_1 ), .B(BIBUF_COREI2C_0_0_SDA_IO_Y), .Y(
        \SDAI_ff_reg_3[0] ));
    CFG4 #( .INIT(16'h1191) )  \fsmmod_ns_0_0_o2_1[3]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(pedetect_net_1), 
        .D(\fsmsta[0]_net_1 ), .Y(\fsmmod_ns_0_0_o2_1[3]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  PRDATA_m6_0_m4 (.A(\sercon[7]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(\sersta[4]_net_1 ), .Y(
        PRDATA_N_9));
    CFG4 #( .INIT(16'hECCC) )  \serdat_write_proc.bsd7_tmp_7s2  (.A(
        un1_PSEL_0), .B(\fsmdet[3]_net_1 ), .C(m3_0), .D(
        CoreAPB3_0_APBmslave0_PSELx), .Y(bsd7_tmp_7_sm0));
    CFG4 #( .INIT(16'h48EA) )  \fsmsta_sync_proc.fsmsta_9_0_o2_6_1[0]  
        (.A(\fsmsta[4]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(
        \fsmsta_9_0_o2_6_1_1[0] ), .D(N_358), .Y(
        \fsmsta_9_0_o2_6_1[0] ));
    CFG3 #( .INIT(8'h02) )  \fsmsta_sync_proc.fsmsta_9_0_a2_0_1[4]  (
        .A(\fsmsta[4]_net_1 ), .B(\fsmdet[3]_net_1 ), .C(framesync24), 
        .Y(\fsmsta_9_0_a2_0_1[4] ));
    CFG4 #( .INIT(16'hDC50) )  \fsmsta_sync_proc.fsmsta_9_0_3[4]  (.A(
        \fsmdet[3]_net_1 ), .B(\fsmsta_9_0_a2_3_1[4] ), .C(N_228), .D(
        N_480_2), .Y(\fsmsta_9_0_3[4] ));
    SLE \SCLI_ff_reg[3]  (.D(N_295_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[3]_net_1 ));
    CFG4 #( .INIT(16'h777F) )  SDAO_int_1_sqmuxa_i (.A(
        SDAO_int_1_sqmuxa_4_net_1), .B(un1_sersta65_1), .C(
        un1_framesync_1), .D(framesync24), .Y(SDAO_int_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'hF4F0) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_6_0  (.A(
        \fsmsta[2]_net_1 ), .B(ack_net_1), .C(N_479), .D(N_542), .Y(
        fsmsta_9_0_372_i_0_o2_6_0));
    CFG2 #( .INIT(4'hD) )  \fsmmod_ns_i_0_o2[4]  (.A(un1_framesync_2), 
        .B(COREI2C_0_0_INT[0]), .Y(N_213));
    CFG2 #( .INIT(4'hD) )  \SCLI_ff_reg_RNO[3]  (.A(\sercon[6]_net_1 ), 
        .B(\SCLI_ff_reg[2]_net_1 ), .Y(N_295_i_0));
    CFG4 #( .INIT(16'hFFFE) )  \fsmsync_sync_proc.un1_fsmsync_2  (.A(
        \fsmsync[2]_net_1 ), .B(\fsmsync[5]_net_1 ), .C(
        \fsmsync[6]_net_1 ), .D(\fsmsync[1]_net_1 ), .Y(un1_fsmsync_2));
    CFG4 #( .INIT(16'hFEFF) )  PCLKint_RNO (.A(
        un14_counter_PRESETN_net_1), .B(un18_counter_PRESETN_net_1), 
        .C(adrcomp12), .D(un1_fsmdet_1_2_net_1), .Y(un1_fsmdet_1_i_0));
    CFG4 #( .INIT(16'hFFDF) )  \fsmmod_ns_0_0_o2[0]  (.A(PCLKint_net_1)
        , .B(N_185), .C(starto_en_net_1), .D(PCLKint_ff_net_1), .Y(
        N_200));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[5]  (.A(
        serdat4), .B(\serdat[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .Y(\serdat_19[5] ));
    CFG4 #( .INIT(16'h4000) )  \SDAO_int_write_proc.un1_framesync_1  (
        .A(\framesync[3]_net_1 ), .B(\framesync[0]_net_1 ), .C(
        \framesync[2]_net_1 ), .D(\framesync[1]_net_1 ), .Y(
        un1_framesync_1));
    CFG4 #( .INIT(16'h0010) )  \PRDATA_0_iv_0_RNO_0[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(\sercon[6]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(sercon_m2_e_2_1));
    CFG4 #( .INIT(16'hF2FA) )  \framesync_write_proc.framesync14_0  (
        .A(sersta77_2), .B(N_394), .C(N_466), .D(N_358), .Y(
        framesync14));
    CFG3 #( .INIT(8'hC8) )  \sercon_write_proc.adrcomp12  (.A(
        \fsmmod[5]_net_1 ), .B(\sercon[4]_net_1 ), .C(
        \fsmmod[0]_net_1 ), .Y(adrcomp12));
    CFG3 #( .INIT(8'hBA) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_1  
        (.A(N_527), .B(framesync24), .C(\fsmsta[3]_net_1 ), .Y(N_395));
    CFG4 #( .INIT(16'hA800) )  un1_ens1_pre_1_sqmuxa_i_a2_1 (.A(N_370), 
        .B(framesync24), .C(un1_framesync24_1), .D(counter_PRESETN_1), 
        .Y(N_514));
    CFG4 #( .INIT(16'h0001) )  \fsmsta_RNO[1]  (.A(
        fsmsta_9_0_372_i_0_3), .B(N_444), .C(fsmsta_9_0_372_i_0_4), .D(
        N_442), .Y(N_1328_i_0));
    CFG4 #( .INIT(16'h8000) )  \serdat_write_proc.serdat4  (.A(
        un12_PSELi), .B(un1_WEn_1), .C(CoreAPB3_0_APBmslave0_PSELx), 
        .D(un4_PRDATA), .Y(serdat4));
    SLE \PCLK_count2[0]  (.D(\PCLK_count2_4[0]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\PCLK_count2[0]_net_1 ));
    SLE \sersta[0]  (.D(\sersta_3[0] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[0]_net_1 ));
    CFG4 #( .INIT(16'h7F20) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_m5  (.A(un1_framesync_1), 
        .B(ack_bit_net_1), .C(un1_sersta65_1), .D(N_1288), .Y(N_1289));
    SLE \PCLK_count1[3]  (.D(\PCLK_count1_4[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[3]_net_1 ));
    SLE \indelay[2]  (.D(\indelay_4[2]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[2]_net_1 ));
    SLE \fsmsync[2]  (.D(N_957_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \sercon_write_proc.sercon_9_0_2[3]  (.A(
        \sercon[6]_net_1 ), .B(N_2_4_tz), .C(\sercon_9_0_0_a0[3] ), .Y(
        \sercon_9_0_0[3] ));
    CFG4 #( .INIT(16'h3777) )  \fsmsync_sync_proc.SCLO_int5_i  (.A(
        un1_fsmsync_2), .B(\sercon[6]_net_1 ), .C(un1_sersta69), .D(
        bsd7_tmp_i_m_1), .Y(SCLO_int5_i_0));
    CFG3 #( .INIT(8'hB8) )  \fsmsta_sync_proc.fsmsta_9_0_m2_ns[2]  (.A(
        \fsmsta_9_0_m2_bm[2] ), .B(framesync24), .C(
        \fsmsta_9_0_m2_am[2] ), .Y(N_226));
    CFG2 #( .INIT(4'h6) )  \sersta_write_proc.sersta_3_0_x2[0]  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[1]_net_1 ), .Y(N_140_i));
    CFG3 #( .INIT(8'hC8) )  \fsmsta_sync_proc.fsmsta_9_0_a2_13[0]  (.A(
        N_496), .B(framesync24), .C(N_497), .Y(N_530));
    CFG4 #( .INIT(16'hE000) )  \fsmdet_RNO[5]  (.A(\fsmdet[2]_net_1 ), 
        .B(\fsmdet[4]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_879_i_0));
    CFG4 #( .INIT(16'h8000) )  \serdat_RNIC4T64[5]  (.A(un12_PSELi), 
        .B(CoreAPB3_0_APBmslave0_PRDATA_m_1[7]), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(\serdat_RNI49U42[5]_net_1 ), 
        .Y(CoreAPB3_0_APBmslave0_PRDATA_m_4));
    CFG4 #( .INIT(16'h7CFC) )  \fsmsta_sync_proc.fsmsta_9_0_o2_4[2]  (
        .A(\fsmsta[0]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \fsmsta[2]_net_1 ), .D(N_367), .Y(N_255));
    SLE \framesync[3]  (.D(\framesync_6[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[3]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \SMBint_filter_proc.SCLI_ff_reg_3[0]  (.A(
        \sercon[6]_net_1 ), .B(BIBUF_COREI2C_0_0_SCL_IO_Y), .Y(
        \SCLI_ff_reg_3[0] ));
    CFG3 #( .INIT(8'h1D) )  \sersta_RNI4IEV[2]  (.A(\sercon[5]_net_1 ), 
        .B(CoreAPB3_0_APBmslave0_PADDR[2]), .C(\sersta[2]_net_1 ), .Y(
        r_N_3_0));
    CFG4 #( .INIT(16'hFFEC) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_3_2  (.A(N_152), .B(
        fsmsta_9_2_342_i_i_o2_3_0), .C(fsmsta_9_2_342_i_i_a2_10_0), .D(
        N_512), .Y(fsmsta_9_2_342_i_i_o2_3_2));
    CFG2 #( .INIT(4'hD) )  \SCLI_ff_reg_RNO[2]  (.A(\sercon[6]_net_1 ), 
        .B(\SCLI_ff_reg[1]_net_1 ), .Y(N_294_i_0));
    CFG4 #( .INIT(16'hFF40) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_10  (.A(
        \fsmsta[4]_net_1 ), .B(framesync24), .C(ack_net_1), .D(
        \fsmsta[3]_net_1 ), .Y(N_152));
    CFG4 #( .INIT(16'h4044) )  \fsmsta_sync_proc.fsmsta_9_0_a2_4_0[0]  
        (.A(ack_net_1), .B(adrcompen_net_1), .C(N_360), .D(
        \fsmsta[2]_net_1 ), .Y(\fsmsta_9_0_a2_4_0[0] ));
    CFG2 #( .INIT(4'hE) )  \fsmmod_ns_i_0_o2_1[2]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_355));
    CFG2 #( .INIT(4'h4) )  \fsmsta_sync_proc.fsmsta_9_0_a2_1_0[4]  (.A(
        \fsmdet[3]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(
        \fsmsta_9_0_a2_2_0[4] ));
    CFG3 #( .INIT(8'h01) )  \adrcomp_write_proc.un1_ack_0_a2_1  (.A(
        \serdat[6]_net_1 ), .B(\serdat[5]_net_1 ), .C(
        \serdat[1]_net_1 ), .Y(un1_ack_1_0));
    CFG4 #( .INIT(16'hF3F2) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_3  (.A(N_151), .B(
        N_356), .C(fsmsta_9_2_342_i_i_o2_3_2), .D(
        fsmsta_9_2_342_i_i_a2_8_0), .Y(N_413));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[0]  (.A(
        serdat4), .B(ack_net_1), .C(CoreAPB3_0_APBmslave0_PWDATA[0]), 
        .Y(\serdat_19[0] ));
    CFG3 #( .INIT(8'h6A) )  \serdat_write_proc.bsd7_10_iv_i_RNO_0  (.A(
        d_N_5_mux), .B(bsd7_N_12_mux), .C(r_N_4_mux), .Y(bsd7_i_m));
    CFG3 #( .INIT(8'hA8) )  \un1_framesync_1_1.CO0  (.A(
        \framesync[0]_net_1 ), .B(nedetect_net_1), .C(un1_framesync_2), 
        .Y(CO0));
    CFG4 #( .INIT(16'h50D8) )  un1_ens1_pre_1_sqmuxa_i_0_1 (.A(
        counter_PRESETN_1), .B(N_380), .C(pedetect_net_1), .D(
        COREI2C_0_0_INT[0]), .Y(un1_ens1_pre_1_sqmuxa_i_0_1_net_1));
    CFG4 #( .INIT(16'h00E0) )  \fsmmod_ns_0_0_a2_0[5]  (.A(N_360), .B(
        N_356), .C(\fsmmod_ns_0_0_a2_0_0[5]_net_1 ), .D(N_372), .Y(
        N_301));
    SLE PCLK_count1_ov (.D(PCLK_count1_ov_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PCLK_count1_ov_net_1));
    CFG3 #( .INIT(8'h80) )  \sersta_write_proc.sersta_3_0_a2_2[1]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[3]_net_1 ), .Y(N_524));
    CFG4 #( .INIT(16'hFD00) )  \sersta_write_proc.sersta_3_0_a2[4]  (
        .A(\fsmsta[1]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(
        \fsmsta[2]_net_1 ), .D(\fsmsta[4]_net_1 ), .Y(N_291));
    CFG3 #( .INIT(8'h08) )  \serdat_write_proc.bsd7_tmp_7_bm  (.A(
        un1_sersta58_0), .B(CoreAPB3_0_APBmslave0_PWDATA[7]), .C(
        \fsmdet[3]_net_1 ), .Y(bsd7_tmp_7_bm));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_RNO[3]  (.A(\sercon[6]_net_1 ), 
        .B(\SDAI_ff_reg[2]_net_1 ), .Y(N_68_i_0));
    CFG4 #( .INIT(16'h0002) )  \fsmsta_sync_proc.fsmsta_9_0_a2_15[0]  
        (.A(ack_net_1), .B(SDAInt_net_1), .C(N_364), .D(N_355), .Y(
        N_496));
    CFG4 #( .INIT(16'hFFFE) )  
        \SCLInt_write_proc.un1_SCLI_ff_reg_i_0_a2  (.A(
        \SCLI_ff_reg[0]_net_1 ), .B(\SCLI_ff_reg[3]_net_1 ), .C(
        \SCLI_ff_reg[2]_net_1 ), .D(\SCLI_ff_reg[1]_net_1 ), .Y(N_262));
    SLE \indelay[1]  (.D(\indelay_4[1]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[1]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \PRDATA_0_iv_0_RNO_0[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(COREI2C_0_0_INT[0]), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(sercon_m2_e_1));
    CFG4 #( .INIT(16'hFAFE) )  \adrcomp_write_proc.un1_sersta64_1  (.A(
        \fsmmod[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmmod[5]_net_1 ), .D(N_360), .Y(un1_sersta64_1));
    CFG4 #( .INIT(16'h0002) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_a2_8_0  (.A(SDAInt_net_1), 
        .B(\fsmsta[3]_net_1 ), .C(\fsmsta[4]_net_1 ), .D(N_358), .Y(
        fsmsta_9_2_342_i_i_a2_8_0));
    CFG4 #( .INIT(16'hF0F4) )  \fsmmod_ns_0_0[1]  (.A(nedetect_net_1), 
        .B(\fsmmod[1]_net_1 ), .C(N_297), .D(N_398), .Y(\fsmmod_ns[1] )
        );
    CFG3 #( .INIT(8'hF2) )  \fsmsync_ns_i_0[6]  (.A(\fsmsync[6]_net_1 )
        , .B(SDAInt_net_1), .C(N_985), .Y(\fsmsync_ns_i_0[6]_net_1 ));
    SLE \serdat[0]  (.D(\serdat_19[0] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(serdat_0));
    CFG4 #( .INIT(16'h7370) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1_1[0]  
        (.A(pedetect_net_1), .B(adrcompen_net_1), .C(N_412), .D(N_543), 
        .Y(\fsmsta_9_0_o2_1_1[0] ));
    CFG4 #( .INIT(16'hFFB0) )  \fsmsta_sync_proc.fsmsta_9_0_1[4]  (.A(
        N_401), .B(N_358), .C(\fsmsta_9_0_a2_0_1[4] ), .D(
        \fsmsta_9_0_0[4] ), .Y(\fsmsta_9_0_1[4] ));
    CFG3 #( .INIT(8'hCD) )  \fsmsta_sync_proc.fsmsta_9_0_m2_am[2]  (.A(
        N_355), .B(N_477), .C(N_367), .Y(\fsmsta_9_0_m2_am[2] ));
    CFG3 #( .INIT(8'h02) )  \fsmsta_sync_proc.fsmsta_9_0_a2_3_1[4]  (
        .A(ack_net_1), .B(\fsmdet[3]_net_1 ), .C(N_359), .Y(
        \fsmsta_9_0_a2_3_1[4] ));
    CFG4 #( .INIT(16'h0222) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_a2_9  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \COREI2C_0_0_SDAO[0] ), .D(\fsmsta[0]_net_1 ), .Y(N_512));
    SLE \framesync[2]  (.D(\framesync_6[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[2]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h2303) )  \SDAO_int_write_proc.un1_sersta58_0  (
        .A(\fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(N_365), .D(
        N_526), .Y(un1_sersta58_0));
    CFG3 #( .INIT(8'h10) )  \framesync_write_proc.framesync14_0_a2_2  
        (.A(\fsmsta[2]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \fsmsta[4]_net_1 ), .Y(N_533));
    CFG3 #( .INIT(8'h80) )  
        \PCLK_counter1_proc.PCLK_count1_4_0_a2_0_1[3]  (.A(
        \PCLK_count1[2]_net_1 ), .B(\PCLK_count1[1]_net_1 ), .C(
        \PCLK_count1[0]_net_1 ), .Y(\PCLK_count1_4_0_a2_0_0[3] ));
    CFG4 #( .INIT(16'h0004) )  \fsmmod_ns_i_0_a2_0_0[2]  (.A(
        \fsmmod[6]_net_1 ), .B(PCLKint_ff_net_1), .C(\fsmmod[1]_net_1 )
        , .D(PCLKint_net_1), .Y(\fsmmod_ns_i_0_a2_0_0[2]_net_1 ));
    CFG3 #( .INIT(8'hFB) )  \sersta_write_proc.sersta_3_0[2]  (.A(
        N_414), .B(COREI2C_0_0_INT[0]), .C(N_543), .Y(\sersta_3[2] ));
    CFG2 #( .INIT(4'h1) )  \fsmsync_ns_0_o3_0_a2_1[0]  (.A(
        \fsmmod[5]_net_1 ), .B(\fsmmod[6]_net_1 ), .Y(N_438_1));
    CFG4 #( .INIT(16'h888B) )  \sercon_RNO[4]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .B(sercon18), .C(adrcomp12), 
        .D(N_418), .Y(N_62_i_0));
    CFG4 #( .INIT(16'h5515) )  \fsmsync_ns_i_a3[5]  (.A(
        \fsmsync[5]_net_1 ), .B(\fsmsync[2]_net_1 ), .C(PCLKint_net_1), 
        .D(PCLKint_ff_net_1), .Y(N_994));
    CFG4 #( .INIT(16'hF2F0) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_0_0  (.A(
        adrcompen_net_1), .B(ack_net_1), .C(N_395), .D(N_227), .Y(
        fsmsta_9_2_342_i_i_o2_0));
    CFG3 #( .INIT(8'h8F) )  adrcomp_2_sqmuxa_i (.A(un1_sercon_1_6), .B(
        un1_sersta64_1), .C(un1_adrcomp14_1), .Y(adrcomp_2_sqmuxa_i_0));
    SLE \sersta[1]  (.D(\sersta_3[1] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[1]_net_1 ));
    CFG4 #( .INIT(16'hAE0C) )  \SDAO_int_write_proc.un1_sersta65_1_1  
        (.A(N_1235), .B(N_549), .C(\fsmsta[4]_net_1 ), .D(N_374), .Y(
        un1_sersta65_1_1));
    SLE \fsmdet[4]  (.D(N_877_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[4]_net_1 ));
    SLE \indelay[0]  (.D(\indelay_4[0]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  un9_PRDATA_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_97_1));
    CFG4 #( .INIT(16'h0200) )  \serdat_write_proc.bsd7_10_iv_1_a0_2  (
        .A(CoreAPB3_0_APBmslave0_PENABLE), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PWRITE), .Y(bsd7_10_iv_1_a0_2));
    CFG2 #( .INIT(4'hB) )  \fsmsta_sync_proc.fsmsta_9_0_o2_7[4]  (.A(
        SDAInt_net_1), .B(\COREI2C_0_0_SDAO[0] ), .Y(N_367));
    SLE \fsmdet[0]  (.D(SCLInt_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[0]_net_1 ));
    SLE \sercon[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[7]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \CoreAPB3_0_APBmslave1_PRDATA_m[0]  (.A(
        GPOUT_reg40_2), .B(TRIG_c[0]), .C(CoreAPB3_0_APBmslave1_PSELx), 
        .D(gpin3_m_2_0[1]), .Y(CoreAPB3_0_APBmslave1_PRDATA_m[0]));
    SLE ack_bit (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), 
        .EN(ack_bit_1_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(ack_bit_net_1));
    CFG3 #( .INIT(8'h10) )  \PRDATA_0_iv_0_RNO[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(sercon_m2_e_2_1), .Y(
        \sercon_m[6] ));
    SLE \fsmsta[2]  (.D(\fsmsta_9[2] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fsmsta[2]_net_1 ));
    CFG4 #( .INIT(16'h0CAE) )  adrcomp_2_sqmuxa_0_1 (.A(sersta77_2), 
        .B(\fsmsta[2]_net_1 ), .C(N_360), .D(N_358), .Y(
        adrcomp_2_sqmuxa_0_1_net_1));
    CFG4 #( .INIT(16'h0008) )  \fsmsta_sync_proc.fsmsta_9_0_a2_7[0]  (
        .A(adrcompen_net_1), .B(ack_net_1), .C(N_360), .D(N_356), .Y(
        N_490));
    CFG3 #( .INIT(8'h01) )  \CoreAPB3_0_APBmslave0_PRDATA_m_1[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[1]), .C(
        CoreAPB3_0_APBmslave0_PADDR[0]), .Y(
        CoreAPB3_0_APBmslave0_PRDATA_m_1[7]));
    CFG4 #( .INIT(16'hF7F3) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_1  (.A(adrcomp_net_1), 
        .B(\sercon[6]_net_1 ), .C(\fsmmod[3]_net_1 ), .D(
        \fsmmod[0]_net_1 ), .Y(SDAO_int_6_0_312_1));
    CFG2 #( .INIT(4'h8) )  \indelay_write_proc.fsmsync_nxt35  (.A(
        \indelay[1]_net_1 ), .B(\indelay[2]_net_1 ), .Y(fsmsync_nxt35));
    SLE \fsmdet[2]  (.D(N_873_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[2]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  \SCLInt_write_proc.SCLInt6_0_a2  (.A(
        \SCLI_ff_reg[0]_net_1 ), .B(\SCLI_ff_reg[3]_net_1 ), .C(
        \SCLI_ff_reg[2]_net_1 ), .D(\SCLI_ff_reg[1]_net_1 ), .Y(
        pedetect_0_sqmuxa_3));
    CFG4 #( .INIT(16'h0E00) )  \fsmdet_RNO[2]  (.A(\fsmdet[0]_net_1 ), 
        .B(\fsmdet[2]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_873_i_0));
    SLE \framesync[1]  (.D(\framesync_6[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[1]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  \serdat_write_proc.bsd7_10_iv_i_RNO  (
        .A(un1_sersta58_0), .B(CoreAPB3_0_APBmslave0_PWDATA[7]), .C(
        COREI2C_0_0_INT[0]), .D(\fsmdet[3]_net_1 ), .Y(
        \PWDATA_i_m_1[7] ));
    CFG4 #( .INIT(16'h0010) )  \sercon_RNI8SHD1[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(\sercon[1]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(sercon_m2_e_3_1));
    SLE \sercon[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(sercon_0));
    CFG4 #( .INIT(16'h0028) )  
        \SDAO_int_write_proc.un1_sersta65_1_2_0_0_a2  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[4]_net_1 ), .D(N_364), .Y(N_460));
    SLE \fsmsync[1]  (.D(N_955_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[1]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \fsmmod_ns_i_0_a2_0[2]  (.A(
        \sercon[5]_net_1 ), .B(COREI2C_0_0_INT[0]), .C(
        \fsmmod_ns_i_0_a2_0_0[2]_net_1 ), .D(
        \fsmmod_ns_i_0_a2_0_2[2]_net_1 ), .Y(N_453));
    CFG3 #( .INIT(8'h40) )  nedetect_RNIGVSG (.A(COREI2C_0_0_INT[0]), 
        .B(un1_sersta58_0), .C(nedetect_net_1), .Y(\serdat_i_m_3_1[7] )
        );
    SLE \fsmmod[0]  (.D(\fsmmod_ns[0] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[0]_net_1 ));
    CFG4 #( .INIT(16'hCECC) )  \SDAO_int_write_proc.un1_sersta65_1_0  
        (.A(N_492), .B(N_460), .C(\fsmsta[1]_net_1 ), .D(N_526), .Y(
        un1_sersta65_1_0));
    CFG4 #( .INIT(16'h0400) )  \fsmsta_sync_proc.fsmsta_9_0_a2_9[2]  (
        .A(N_367), .B(\fsmsta[0]_net_1 ), .C(N_364), .D(N_492), .Y(
        N_476));
    CFG4 #( .INIT(16'hECCC) )  \PRDATA_0_iv_0[3]  (.A(N_97_1), .B(
        \sercon_m[3] ), .C(\sersta[0]_net_1 ), .D(un9_PRDATA_1_net_1), 
        .Y(\PRDATA_0_iv_0[3]_net_1 ));
    SLE \fsmmod[6]  (.D(N_1016_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[6]_net_1 ));
    CFG4 #( .INIT(16'hFF10) )  \fsmmod_ns_i_0_o2[6]  (.A(N_360), .B(
        N_356), .C(pedetect_net_1), .D(N_372), .Y(N_398));
    SLE \sercon[4]  (.D(N_62_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sercon[4]_net_1 ));
    CFG3 #( .INIT(8'h09) )  un1_ens1_pre_1_sqmuxa_i_o2_0 (.A(
        \framesync[3]_net_1 ), .B(\framesync[0]_net_1 ), .C(N_1028_2), 
        .Y(N_380));
    CFG4 #( .INIT(16'h2303) )  \fsmsta_sync_proc.fsmsta_9_0_1_1[0]  (
        .A(un1_framesync24), .B(N_527), .C(counter_PRESETN_1), .D(
        N_370), .Y(\fsmsta_9_0_1_1[0] ));
    SLE SCLO_int (.D(SCLO_int5_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \COREI2C_0_0_SCLO[0] ));
    SLE \fsmmod[2]  (.D(N_1010_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[2]_net_1 ));
    SLE \sersta[3]  (.D(\sersta_3[3] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[3]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \fsmmod_ns_i_0_a2_1[2]  (.A(
        \fsmmod[1]_net_1 ), .B(N_213), .C(\sercon[4]_net_1 ), .D(
        \fsmmod[6]_net_1 ), .Y(N_455));
    SLE \fsmsync[6]  (.D(N_965_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[6]_net_1 ));
    SLE \SDAI_ff_reg[2]  (.D(N_66_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[2]_net_1 ));
    SLE \fsmsync[0]  (.D(\fsmsync_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[0]_net_1 ));
    CFG4 #( .INIT(16'hA2A0) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_4  (.A(framesync24), 
        .B(N_360), .C(pedetect_net_1), .D(\fsmsta[2]_net_1 ), .Y(N_227)
        );
    SLE \PCLK_count1[0]  (.D(N_340_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[0]_net_1 ));
    CFG4 #( .INIT(16'hFFCA) )  \sercon_write_proc.sercon_9_0[3]  (.A(
        COREI2C_0_0_INT[0]), .B(CoreAPB3_0_APBmslave0_PWDATA[3]), .C(
        sercon18), .D(\sercon_9_0_0[3] ), .Y(\sercon_9[3] ));
    CFG3 #( .INIT(8'hEF) )  \fsmmod_ns_0_0_o2_2[3]  (.A(
        \sercon[4]_net_1 ), .B(COREI2C_0_0_INT[0]), .C(
        \sercon[5]_net_1 ), .Y(N_185));
    SLE \fsmsta[0]  (.D(\fsmsta_9[0] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fsmsta[0]_net_1 ));
    SLE \serdat[3]  (.D(\serdat_19[3] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \sercon_write_proc.un1_PSEL_0  (.A(
        CoreAPB3_0_APBmslave0_PENABLE), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .Y(un1_WEn_1));
    SLE nedetect (.D(nedetect_0_sqmuxa), .CLK(GL0_INST), .EN(
        pedetect_0_sqmuxa_3), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(nedetect_net_1));
    CFG4 #( .INIT(16'h0400) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_18  (.A(
        \fsmsta_9_0_o2_3_0[2] ), .B(\fsmsta[4]_net_1 ), .C(N_356), .D(
        N_358), .Y(N_509));
    CFG4 #( .INIT(16'hECCC) )  \fsmmod_ns_0_0_0[0]  (.A(
        \fsmmod[5]_net_1 ), .B(N_548), .C(sclscl_net_1), .D(
        pedetect_net_1), .Y(\fsmmod_ns_0_0_0[0]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \sersta_write_proc.sersta_3_0_a2_4[3]  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \fsmsta[2]_net_1 ), .Y(N_549));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.bsd7_tmp_7_ns  (.A(
        bsd7_tmp_7_sm0), .B(bsd7_tmp_7_am), .C(bsd7_tmp_7_bm), .Y(
        bsd7_tmp_7));
    CFG3 #( .INIT(8'h08) )  un1_ens1_pre_1_sqmuxa_i_a2_2 (.A(
        \fsmmod[4]_net_1 ), .B(PCLKint_ff_net_1), .C(PCLKint_net_1), 
        .Y(N_527));
    CFG4 #( .INIT(16'hCECC) )  \fsmsta_sync_proc.fsmsta_9_0_o2_3_0[0]  
        (.A(\fsmsta[0]_net_1 ), .B(N_527), .C(framesync24), .D(N_384), 
        .Y(\fsmsta_9_0_o2_3_0[0] ));
    CFG4 #( .INIT(16'hFFEA) )  adrcompen_2_sqmuxa_i (.A(adrcomp12), .B(
        framesync24), .C(nedetect_net_1), .D(\fsmdet[3]_net_1 ), .Y(
        adrcompen_2_sqmuxa_i_0));
    CFG2 #( .INIT(4'h4) )  \sersta_write_proc.sersta_3_0_a2_2[3]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_531));
    CFG4 #( .INIT(16'h4000) )  \serdat_write_proc.bsd7_10_iv_i_RNO_2  
        (.A(bsd7_net_1), .B(un1_sersta58_0), .C(un1_WEn_1), .D(
        bsd7_m6_3), .Y(bsd7_N_12_mux));
    CFG3 #( .INIT(8'hF7) )  \sersta_write_proc.sersta_3_0[0]  (.A(
        N_224), .B(COREI2C_0_0_INT[0]), .C(N_526), .Y(\sersta_3[0] ));
    CFG1 #( .INIT(2'h1) )  SCLO_int_RNI12J6 (.A(\COREI2C_0_0_SCLO[0] ), 
        .Y(COREI2C_0_0_SCLO_i[0]));
    CFG4 #( .INIT(16'h3ACA) )  
        \framesync_write_proc.framesync_6_enl[1]  (.A(
        \fsmdet[3]_net_1 ), .B(\framesync[1]_net_1 ), .C(
        framesync_6_e2), .D(CO0), .Y(\framesync_6[1] ));
    CFG4 #( .INIT(16'hA8A0) )  \CoreAPB3_0_APBmslave1_PRDATA_m[1]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(GPOUT_reg[1]), .C(gpin3_m[1]), 
        .D(GPOUT_reg40), .Y(CoreAPB3_0_APBmslave1_PRDATA_m[1]));
    CFG3 #( .INIT(8'hFE) )  \serdat_write_proc.un1_sersta65  (.A(
        un1_sersta65_1), .B(\fsmdet[3]_net_1 ), .C(un1_sersta58_0), .Y(
        un1_sersta65));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_RNO[1]  (.A(\sercon[6]_net_1 ), 
        .B(\SDAI_ff_reg[0]_net_1 ), .Y(N_64_i_0));
    CFG2 #( .INIT(4'hE) )  \fsmsync_ns_i_o3[3]  (.A(N_994), .B(
        COREI2C_0_0_INT[0]), .Y(N_973));
    CFG2 #( .INIT(4'hE) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_1  
        (.A(fsmsta_9_0_372_i_0_o2_1_4), .B(N_509), .Y(N_404));
    CFG4 #( .INIT(16'hFFFB) )  \fsmsta_sync_proc.fsmsta_9_0_o2_9[0]  (
        .A(SDAInt_net_1), .B(\COREI2C_0_0_SDAO[0] ), .C(N_365), .D(
        \fsmsta[3]_net_1 ), .Y(N_384));
    CFG2 #( .INIT(4'h8) )  \CoreAPB3_0_APBmslave0_PRDATA_m_0[1]  (.A(
        CoreAPB3_0_APBmslave0_PSELx), .B(un12_PSELi), .Y(
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]));
    CFG4 #( .INIT(16'hCCEC) )  \serdat_write_proc.ack_10_u_xx  (.A(
        COREI2C_0_0_INT[0]), .B(ack_net_1), .C(un1_sersta58_0), .D(
        \fsmdet[3]_net_1 ), .Y(ack_10_u_xx));
    CFG4 #( .INIT(16'hFFB3) )  \sersta_write_proc.sersta_3_0_1[3]  (.A(
        N_416), .B(COREI2C_0_0_INT[0]), .C(N_492), .D(N_531), .Y(
        \sersta_3_0_1[3] ));
    CFG4 #( .INIT(16'h0013) )  \PCLK_count1_RNO[0]  (.A(
        \PCLK_count1[3]_net_1 ), .B(\PCLK_count1[0]_net_1 ), .C(N_155), 
        .D(counter_PRESETN_net_1), .Y(N_340_i_0));
    CFG4 #( .INIT(16'h0405) )  SDAO_int_1_sqmuxa_1 (.A(
        \fsmmod[6]_net_1 ), .B(adrcomp_net_1), .C(\fsmmod[4]_net_1 ), 
        .D(\fsmmod[0]_net_1 ), .Y(SDAO_int_1_sqmuxa_1_net_1));
    SLE \fsmsta[1]  (.D(N_1328_i_0), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\fsmsta[1]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \adrcomp_write_proc.un1_sercon_1_5  (.A(
        un1_framesync_1), .B(N_244), .Y(un1_sercon_1_5));
    CFG4 #( .INIT(16'hFFFB) )  \sersta_write_proc.sersta_3_0[4]  (.A(
        sersta77_2), .B(COREI2C_0_0_INT[0]), .C(N_292), .D(N_291), .Y(
        \sersta_3[4] ));
    CFG4 #( .INIT(16'hFF2A) )  \serdat_write_proc.bsd7_tmp_7_am  (.A(
        \serdat_i_m_3_1[7] ), .B(un1_PSEL_0), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(\serdat_i_m_3_0_0[7] ), .Y(
        bsd7_tmp_7_am));
    CFG4 #( .INIT(16'h0010) )  un1_fsmdet_1_2 (.A(\fsmdet[5]_net_1 ), 
        .B(PCLK_count2_ov_net_1), .C(N_827), .D(\fsmdet[3]_net_1 ), .Y(
        un1_fsmdet_1_2_net_1));
    SLE \SDAI_ff_reg[3]  (.D(N_68_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[3]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \fsmsta_sync_proc.fsmsta_9_0_a2_3_2[4]  (
        .A(\fsmsta[0]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(N_356), .Y(
        N_480_2));
    SLE \framesync[0]  (.D(\framesync_6[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[0]_net_1 ));
    SLE bsd7_tmp (.D(bsd7_tmp_7), .CLK(GL0_INST), .EN(
        \sercon[6]_net_1 ), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(bsd7_tmp_net_1));
    SLE \fsmdet[3]  (.D(N_875_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[3]_net_1 ));
    CFG3 #( .INIT(8'h01) )  un1_counter_PRESETN_i_a2 (.A(
        \fsmsync[1]_net_1 ), .B(\fsmsync[5]_net_1 ), .C(
        \fsmsync[4]_net_1 ), .Y(N_827));
    CFG4 #( .INIT(16'hECCC) )  \PRDATA_0_iv_0[4]  (.A(N_97_1), .B(
        \sercon_m[4] ), .C(\sersta[1]_net_1 ), .D(un9_PRDATA_1_net_1), 
        .Y(\PRDATA_0_iv_0[4]_net_1 ));
    CFG4 #( .INIT(16'h0051) )  \serdat_write_proc.bsd7_10_iv_1_a1  (.A(
        bsd7_tmp_i_m_1_0), .B(\serdat_i_m_3_1[7] ), .C(
        \serdat[7]_net_1 ), .D(\fsmdet[3]_net_1 ), .Y(bsd7_10_iv_1_a1));
    SLE PCLKint_ff (.D(PCLKint_ff_3), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PCLKint_ff_net_1));
    SLE \serdat[6]  (.D(\serdat_19[6] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[6]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \fsmsta_sync_proc.fsmsta_9_0_a2_7[2]  (
        .A(\fsmsta[1]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(N_526), 
        .D(\fsmsta[4]_net_1 ), .Y(N_474));
    CFG1 #( .INIT(2'h1) )  \fsmdet_RNO[0]  (.A(SCLInt_net_1), .Y(
        SCLInt_i_0));
    CFG4 #( .INIT(16'h0001) )  \fsmmod_RNO[2]  (.A(N_452), .B(N_398), 
        .C(N_455), .D(N_453), .Y(N_1010_i_0));
    CFG4 #( .INIT(16'hFFFE) )  
        \adrcomp_write_proc.un1_sercon_1_8_i_o2  (.A(\serdat[4]_net_1 )
        , .B(\serdat[3]_net_1 ), .C(serdat_2), .D(serdat_0), .Y(N_244));
    CFG4 #( .INIT(16'hBAFF) )  \fsmmod_ns_0_0_o2[3]  (.A(N_355), .B(
        framesync24), .C(\fsmsta[2]_net_1 ), .D(
        \fsmmod_ns_0_0_o2_1[3]_net_1 ), .Y(N_162));
    CFG3 #( .INIT(8'hB7) )  \fsmmod_ns_i_0_o2_3[6]  (.A(PCLKint_net_1), 
        .B(SCLInt_net_1), .C(PCLKint_ff_net_1), .Y(N_407));
    CFG3 #( .INIT(8'h3B) )  starto_en_1_sqmuxa_i_0 (.A(PCLKint_net_1), 
        .B(N_344), .C(PCLKint_ff_net_1), .Y(
        starto_en_1_sqmuxa_i_0_net_1));
    CFG4 #( .INIT(16'h1333) )  
        \sercon_write_proc.sercon_9_0_0_a1_tz_0[3]  (.A(framesync24), 
        .B(N_548), .C(pedetect_net_1), .D(N_370), .Y(
        \sercon_9_0_0_a1_tz_0[3] ));
    CFG4 #( .INIT(16'h000B) )  \fsmmod_RNO[6]  (.A(\fsmmod[3]_net_1 ), 
        .B(nedetect_net_1), .C(N_317), .D(N_398), .Y(N_1016_i_0));
    SLE bsd7 (.D(bsd7_10_iv_i_0), .CLK(GL0_INST), .EN(
        \sercon[6]_net_1 ), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(bsd7_net_1));
    SLE PCLKint (.D(PCLKint_4), .CLK(GL0_INST), .EN(un1_fsmdet_1_i_0), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PCLKint_net_1));
    CFG4 #( .INIT(16'hFF0D) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_i_0  
        (.A(adrcomp_net_1), .B(un1_framesync24), .C(N_221), .D(N_527), 
        .Y(fsmsta_9_2_342_i_i_0));
    SLE \PCLK_count1[1]  (.D(N_341_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[1]_net_1 ));
    SLE \serdat[5]  (.D(\serdat_19[5] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[5]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \sercon_write_proc.sercon_9_0_a2_0_1[3]  (
        .A(adrcomp_net_1), .B(counter_PRESETN_1), .C(N_380), .Y(
        \sercon_9_0_a2_0_1[3] ));
    CFG4 #( .INIT(16'hECCC) )  \fsmsync_ns_0[0]  (.A(N_972), .B(
        \fsmsync_ns_0_1[0]_net_1 ), .C(\fsmsync[0]_net_1 ), .D(
        SCLInt_net_1), .Y(\fsmsync_ns[0] ));
    CFG3 #( .INIT(8'h10) )  \fsmsta_sync_proc.fsmsta_9_0_a2_8_0[2]  (
        .A(SDAInt_net_1), .B(\fsmsta[2]_net_1 ), .C(ack_net_1), .Y(
        \fsmsta_9_0_a2_8_0[2] ));
    CFG4 #( .INIT(16'h0010) )  \serdat_write_proc.bsd7_10_iv_1_a0_3  (
        .A(CoreAPB3_0_APBmslave0_PADDR[7]), .B(\fsmdet[3]_net_1 ), .C(
        bsd7_10_iv_1_a0_2), .D(CoreAPB3_0_APBmslave0_PADDR[8]), .Y(
        bsd7_10_iv_1_a0_3));
    CFG3 #( .INIT(8'hCE) )  \fsmsta_sync_proc.fsmsta_9_0[2]  (.A(N_226)
        , .B(N_527), .C(counter_PRESETN_1), .Y(\fsmsta_9[2] ));
    CFG2 #( .INIT(4'h7) )  \sersta_write_proc.sersta_3_0_o2[1]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_361));
    CFG4 #( .INIT(16'h5F1B) )  \fsmmod_ns_i_0_0[4]  (.A(
        \fsmmod[2]_net_1 ), .B(\fsmmod[4]_net_1 ), .C(
        \sercon[4]_net_1 ), .D(N_547), .Y(\fsmmod_ns_i_0_0[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_a2_10_0  (.A(SDAInt_net_1)
        , .B(\fsmsta[1]_net_1 ), .C(\fsmsta[2]_net_1 ), .Y(
        fsmsta_9_2_342_i_i_a2_10_0));
    CFG4 #( .INIT(16'h8000) )  \sercon_write_proc.sercon_9_0_0_a0[3]  
        (.A(un1_PRDATA), .B(CoreAPB3_0_APBmslave0_PSELx), .C(
        un12_PSELi_0), .D(bsd7_10_iv_1_a0_2), .Y(\sercon_9_0_0_a0[3] ));
    CFG4 #( .INIT(16'h0405) )  \fsmsync_RNO[4]  (.A(SCLInt_net_1), .B(
        \fsmsync[4]_net_1 ), .C(N_985), .D(N_980), .Y(N_961_i_0));
    CFG3 #( .INIT(8'h7F) )  \fsmsta_sync_proc.fsmsta_9_0_o2[4]  (.A(
        adrcomp_net_1), .B(pedetect_net_1), .C(adrcompen_net_1), .Y(
        N_129));
    CFG3 #( .INIT(8'h20) )  \fsmsta_sync_proc.fsmsta_9_0_a2_2_2[4]  (
        .A(\fsmsta_9_0_a2_2_0[4] ), .B(N_358), .C(
        \COREI2C_0_0_SDAO[0] ), .Y(\fsmsta_9_0_a2_2_2[4] ));
    CFG4 #( .INIT(16'hFFEF) )  \fsmmod_ns_0_0_o2_0[5]  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(\fsmsta[4]_net_1 ), .Y(N_360));
    SLE \SDAI_ff_reg[0]  (.D(\SDAI_ff_reg_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \fsmsync_RNO[5]  (.A(COREI2C_0_0_INT[0]), 
        .B(N_994), .C(N_985), .Y(N_963_i_0));
    CFG4 #( .INIT(16'hC080) )  
        \serdat_write_proc.un4_PRDATA_1_RNIUOL64  (.A(\sercon_m[1] ), 
        .B(un12_PSELi), .C(CoreAPB3_0_APBmslave0_PSELx), .D(
        \serdat_m[1] ), .Y(CoreAPB3_0_APBmslave0_PRDATA_m_0_d0));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[6]  (.A(
        serdat4), .B(\serdat[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .Y(\serdat_19[6] ));
    CFG4 #( .INIT(16'h1000) )  \fsmmod_ns_0_0_a2_1_0[3]  (.A(
        PCLKint_net_1), .B(N_372), .C(\fsmmod[2]_net_1 ), .D(
        PCLKint_ff_net_1), .Y(\fsmmod_ns_0_0_a2_1[3] ));
    SLE adrcomp (.D(un1_adrcomp14_1), .CLK(GL0_INST), .EN(
        adrcomp_2_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(adrcomp_net_1));
    CFG4 #( .INIT(16'hFFF8) )  serdat_1_sqmuxa_1_RNIL62J1 (.A(
        \sercon[6]_net_1 ), .B(serdat_2_sqmuxa_out), .C(
        serdat_1_sqmuxa_1_net_1), .D(bsd7_10_iv_1_a0_2_RNI6O401), .Y(
        un1_N_9_mux_i_0));
    CFG4 #( .INIT(16'h0010) )  
        \sercon_write_proc.sercon_9_0_0_a1_tz[3]  (.A(N_514), .B(N_443)
        , .C(\sercon_9_0_0_a1_tz_0[3] ), .D(\sercon_9_0_a2_0_1[3] ), 
        .Y(N_2_4_tz));
    CFG4 #( .INIT(16'h0004) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_a5_0  (.A(
        \fsmmod[1]_net_1 ), .B(N_359), .C(\fsmmod[4]_net_1 ), .D(
        \fsmmod[6]_net_1 ), .Y(SDAO_int_6_0_312_a5_0));
    CFG2 #( .INIT(4'hE) )  \PCLKint_write_proc.PCLKint_ff_3  (.A(
        counter_PRESETN_net_1), .B(PCLKint_net_1), .Y(PCLKint_ff_3));
    CFG3 #( .INIT(8'h0D) )  \serdat_write_proc.bsd7_10_iv_i_RNO_4  (.A(
        nedetect_net_1), .B(COREI2C_0_0_INT[0]), .C(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(bsd7_m6_0));
    SLE adrcompen (.D(un1_adrcomp14_net_1), .CLK(GL0_INST), .EN(
        adrcompen_2_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(adrcompen_net_1));
    CFG4 #( .INIT(16'hCCCE) )  \fsmsync_ns_i_0[3]  (.A(fsmsync_nxt35), 
        .B(N_985), .C(\fsmsync[2]_net_1 ), .D(\fsmsync[5]_net_1 ), .Y(
        \fsmsync_ns_i_0[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \sersta_write_proc.sersta_3_0_m2[0]  (.A(
        \fsmsta[0]_net_1 ), .B(N_140_i), .C(N_361), .Y(N_224));
    SLE \SDAI_ff_reg[1]  (.D(N_64_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hF7F0) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2  (.A(adrcompen_net_1), 
        .B(pedetect_net_1), .C(fsmsta_9_2_342_i_i_o2_0), .D(N_413), .Y(
        N_117));
    CFG2 #( .INIT(4'h4) )  \sersta_write_proc.sersta_3_0_a2_0[3]  (.A(
        N_361), .B(N_394), .Y(N_289));
    CFG3 #( .INIT(8'h08) )  \SDAO_int_write_proc.SDAO_int6  (.A(
        \framesync[0]_net_1 ), .B(nedetect_net_1), .C(
        \framesync[3]_net_1 ), .Y(SDAO_int6));
    CFG4 #( .INIT(16'h11B3) )  \fsmsta_sync_proc.fsmsta_9_0_1[0]  (.A(
        \fsmdet[3]_net_1 ), .B(\fsmsta_9_0_1_1[0] ), .C(
        \fsmmod[6]_net_1 ), .D(\fsmmod[1]_net_1 ), .Y(
        \fsmsta_9_0_1[0] ));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[1]  (.A(
        serdat4), .B(serdat_0), .C(CoreAPB3_0_APBmslave0_PWDATA[1]), 
        .Y(\serdat_19[1] ));
    CFG4 #( .INIT(16'h2000) )  PCLK_count2_ov_0_sqmuxa (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN_net_1), .C(
        \PCLK_count2[1]_net_1 ), .D(\PCLK_count2[0]_net_1 ), .Y(
        PCLK_count2_ov_0_sqmuxa_net_1));
    CFG4 #( .INIT(16'h5054) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_11  (.A(N_129), .B(
        \fsmsta[2]_net_1 ), .C(fsmsta_9_0_372_i_0_o2_12_1), .D(N_360), 
        .Y(N_551));
    SLE \fsmdet[6]  (.D(N_881_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[6]_net_1 ));
    CFG4 #( .INIT(16'hF4F0) )  \serdat_write_proc.ack_10_u_yy  (.A(
        \fsmdet[3]_net_1 ), .B(un1_sersta58_0), .C(SDAInt_net_1), .D(
        COREI2C_0_0_INT[0]), .Y(ack_10_u_yy));
    CFG3 #( .INIT(8'h7F) )  \fsmsync_ns_i_o3[4]  (.A(
        \indelay[1]_net_1 ), .B(\indelay[2]_net_1 ), .C(
        \fsmsync[3]_net_1 ), .Y(N_980));
    CFG4 #( .INIT(16'h0004) )  \serdat_write_proc.bsd7_10_iv_i_RNO_1  
        (.A(COREI2C_0_0_INT[0]), .B(un1_sersta58_0), .C(bsd7_net_1), 
        .D(nedetect_net_1), .Y(d_N_5_mux));
    CFG4 #( .INIT(16'h0102) )  \PCLK_count1_RNO[1]  (.A(
        \PCLK_count1[0]_net_1 ), .B(\PCLK_count1[3]_net_1 ), .C(
        counter_PRESETN_net_1), .D(\PCLK_count1[1]_net_1 ), .Y(
        N_341_i_0));
    CFG4 #( .INIT(16'hFF04) )  \fsmmod_ns_0_0_0[5]  (.A(pedetect_net_1)
        , .B(\fsmmod[5]_net_1 ), .C(N_372), .D(N_301), .Y(
        \fsmmod_ns_0_0_0[5]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \fsmmod_ns_i_0_a2_1[4]  (.A(PCLKint_net_1), 
        .B(SCLInt_net_1), .C(PCLKint_ff_net_1), .Y(N_547));
    CFG4 #( .INIT(16'h8000) )  ack_bit_1_sqmuxa (.A(serdat48), .B(
        sercon18), .C(COREI2C_0_0_INT[0]), .D(\sercon[6]_net_1 ), .Y(
        ack_bit_1_sqmuxa_net_1));
    CFG3 #( .INIT(8'hFE) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1_4[2]  (
        .A(N_476), .B(\fsmsta_9_0_o2_1_0[2] ), .C(N_471), .Y(
        \fsmsta_9_0_o2_1_3[2] ));
    CFG3 #( .INIT(8'h01) )  \sercon_write_proc.un1_PRDATA_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(un1_WEn_0));
    CFG2 #( .INIT(4'h6) )  \sersta_write_proc.sersta_3_0_o2_0[1]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_374));
    CFG2 #( .INIT(4'h4) )  \serdat_write_proc.un4_PRDATA_1  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(un4_PRDATA_1));
    CFG3 #( .INIT(8'hFE) )  \SDAO_int_write_proc.un1_sersta65_1  (.A(
        un1_sersta65_1_0), .B(N_1236), .C(un1_sersta65_1_1), .Y(
        un1_sersta65_1));
    CFG4 #( .INIT(16'h0002) )  \SDAO_int_write_proc.framesync24  (.A(
        \framesync[3]_net_1 ), .B(\framesync[0]_net_1 ), .C(
        \framesync[2]_net_1 ), .D(\framesync[1]_net_1 ), .Y(
        framesync24));
    CFG4 #( .INIT(16'h0103) )  adrcomp_2_sqmuxa_0 (.A(
        COREI2C_0_0_INT[0]), .B(adrcomp12), .C(adrcomp7_0_0), .D(
        adrcomp_2_sqmuxa_0_1_net_1), .Y(un1_adrcomp14_1));
    CFG4 #( .INIT(16'h0040) )  serdat_2_sqmuxa_s (.A(
        COREI2C_0_0_INT[0]), .B(pedetect_net_1), .C(un1_sersta58_0), 
        .D(\fsmdet[3]_net_1 ), .Y(serdat_2_sqmuxa_out));
    SLE \sersta[4]  (.D(\sersta_3[4] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[4]_net_1 ));
    SLE SCLInt (.D(\SCLI_ff_reg[3]_net_1 ), .CLK(GL0_INST), .EN(
        un1_SCLInt5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        SCLInt_net_1));
    CFG4 #( .INIT(16'h0001) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_0_0  (.A(
        \fsmdet[3]_net_1 ), .B(N_359), .C(\fsmdet[5]_net_1 ), .D(
        pedetect_net_1), .Y(fsmsta_9_0_372_i_0_a2_0_0));
    CFG3 #( .INIT(8'h08) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_21  (.A(framesync24), 
        .B(SDAInt_net_1), .C(N_355), .Y(N_542));
    CFG3 #( .INIT(8'h37) )  \framesync_write_proc.un1_sersta58  (.A(
        N_355), .B(\sercon[5]_net_1 ), .C(N_364), .Y(un1_sersta58));
    CFG4 #( .INIT(16'hF1F0) )  \fsmsync_ns_i_0[2]  (.A(
        \fsmsync[0]_net_1 ), .B(\fsmsync[1]_net_1 ), .C(N_985), .D(
        N_979), .Y(\fsmsync_ns_i_0[2]_net_1 ));
    SLE PCLK_count2_ov (.D(PCLK_count2_ov_0_sqmuxa_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PCLK_count2_ov_net_1));
    CFG2 #( .INIT(4'h4) )  un1_adrcomp14 (.A(adrcomp12), .B(
        \fsmdet[3]_net_1 ), .Y(un1_adrcomp14_net_1));
    CFG4 #( .INIT(16'hE000) )  \un1_framesync_1_1.CO1  (.A(
        nedetect_net_1), .B(un1_framesync_2), .C(\framesync[1]_net_1 ), 
        .D(\framesync[0]_net_1 ), .Y(CO1));
    CFG4 #( .INIT(16'h1303) )  \fsmsync_RNO[2]  (.A(N_972), .B(
        \fsmsync_ns_i_0[2]_net_1 ), .C(\fsmsync[0]_net_1 ), .D(
        SCLInt_net_1), .Y(N_957_i_0));
    SLE \sercon[3]  (.D(\sercon_9[3] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        COREI2C_0_0_INT[0]));
    CFG4 #( .INIT(16'hF8F0) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_1_3  (.A(framesync24), 
        .B(\COREI2C_0_0_SDAO[0] ), .C(fsmsta_9_0_372_i_0_o2_1_1), .D(
        N_1236), .Y(fsmsta_9_0_372_i_0_o2_1_3));
    SLE \fsmmod[5]  (.D(\fsmmod_ns[5] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[5]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_14  (.A(
        \fsmsta[0]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(N_356), .D(
        N_355), .Y(N_479));
    CFG3 #( .INIT(8'h40) )  \PCLK_counter1_proc.PCLK_count1_ov_3  (.A(
        counter_PRESETN_net_1), .B(\PCLK_count1[3]_net_1 ), .C(N_220), 
        .Y(PCLK_count1_ov_3));
    CFG3 #( .INIT(8'h10) )  un18_counter_PRESETN (.A(SCLInt_net_1), .B(
        \fsmmod[5]_net_1 ), .C(busfree_net_1), .Y(
        un18_counter_PRESETN_net_1));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[7]  (.A(
        serdat4), .B(\serdat[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .Y(\serdat_19[7] ));
    CFG4 #( .INIT(16'h10FF) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_i_o2_3_0  (.A(
        \COREI2C_0_0_SDAO[0] ), .B(\fsmsta[0]_net_1 ), .C(N_531), .D(
        N_361), .Y(fsmsta_9_2_342_i_i_o2_3_0));
    SLE \fsmdet[5]  (.D(N_879_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[5]_net_1 ));
    SLE \fsmmod[1]  (.D(\fsmmod_ns[1] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[1]_net_1 ));
    CFG4 #( .INIT(16'hDC00) )  \fsmdet_RNO[4]  (.A(SDAInt_net_1), .B(
        \fsmdet[3]_net_1 ), .C(\fsmdet[4]_net_1 ), .D(SCLInt_net_1), 
        .Y(N_877_i_0));
    CFG4 #( .INIT(16'hE000) )  \fsmdet_RNO[1]  (.A(\fsmdet[0]_net_1 ), 
        .B(\fsmdet[1]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_871_i_0));
    CFG2 #( .INIT(4'hB) )  \sersta_write_proc.sersta_3_0_o2_1[1]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_393));
    SLE \fsmsync[4]  (.D(N_961_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[4]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \PRDATA_0_iv_0_RNO[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(sercon_m2_e_0_1), .Y(
        \sercon_m[4] ));
    CFG2 #( .INIT(4'hD) )  sclscl_1_sqmuxa_i (.A(\fsmmod[5]_net_1 ), 
        .B(pedetect_net_1), .Y(sclscl_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'hFFFE) )  counter_PRESETN (.A(
        un18_counter_PRESETN_net_1), .B(un14_counter_PRESETN_net_1), 
        .C(counter_PRESETN_0_net_1), .D(adrcomp12), .Y(
        counter_PRESETN_net_1));
    CFG2 #( .INIT(4'hE) )  \fsmmod_ns_i_o4_2[4]  (.A(
        \framesync[1]_net_1 ), .B(\framesync[2]_net_1 ), .Y(N_1028_2));
    CFG4 #( .INIT(16'h0080) )  
        \fsmsync_sync_proc.un1_sersta69_1_a5_1_0_a2  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(\fsmsta[4]_net_1 ), .Y(N_1236));
    CFG4 #( .INIT(16'h1011) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_3_1  (.A(
        fsmsta_9_0_372_i_0_o2_6_0), .B(N_480), .C(framesync24), .D(
        N_554), .Y(fsmsta_9_0_372_i_0_a2_3_1));
    SLE \sercon[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  SCLInt_RNIEO25 (.A(COREI2C_0_0_INT[0]), .B(
        SCLInt_net_1), .Y(bsd7_tmp_i_m_1));
    CFG4 #( .INIT(16'h008A) )  \fsmsync_ns_i_a3[3]  (.A(
        \sercon[4]_net_1 ), .B(un1_framesync_2), .C(\fsmsync[2]_net_1 )
        , .D(\fsmsync[3]_net_1 ), .Y(N_990));
    CFG2 #( .INIT(4'h2) )  \sersta_write_proc.sersta_3_0_a2[0]  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_526));
    CFG4 #( .INIT(16'h4532) )  
        \fsmsta_sync_proc.fsmsta_9_0_o2_6_1_1[0]  (.A(
        \fsmsta[3]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(N_365), .D(
        \fsmsta[4]_net_1 ), .Y(\fsmsta_9_0_o2_6_1_1[0] ));
    CFG4 #( .INIT(16'h4000) )  \serdat_write_proc.bsd7_tmp_7_sn.m3_0  
        (.A(\fsmdet[3]_net_1 ), .B(COREI2C_0_0_INT[0]), .C(un4_PRDATA), 
        .D(un1_sersta58_0), .Y(m3_0));
    CFG4 #( .INIT(16'h13FF) )  \framesync_write_proc.framesync_6[0]  (
        .A(framesync14), .B(framesync10), .C(un1_framesync_2), .D(
        framesync_6_e2_1), .Y(\framesync_6_m2[3] ));
    CFG4 #( .INIT(16'hA020) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_17  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \fsmsta[4]_net_1 ), .D(\fsmsta[2]_net_1 ), .Y(N_507));
    CFG4 #( .INIT(16'hDCCC) )  \adrcomp_write_proc.adrcomp7_0_0  (.A(
        N_394), .B(counter_PRESETN_1), .C(COREI2C_0_0_INT[0]), .D(
        \fsmsta[4]_net_1 ), .Y(adrcomp7_0_0));
    CFG2 #( .INIT(4'hD) )  \SCLI_ff_reg_RNO[1]  (.A(\sercon[6]_net_1 ), 
        .B(\SCLI_ff_reg[0]_net_1 ), .Y(N_293_i_0));
    CFG4 #( .INIT(16'hF080) )  \PRDATA_0_iv_0_RNI2NIF1[6]  (.A(
        un4_PRDATA), .B(\serdat[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]), .D(
        \PRDATA_0_iv_0[6]_net_1 ), .Y(CoreAPB3_0_APBmslave0_PRDATA_m_5)
        );
    CFG4 #( .INIT(16'hD000) )  serdat_1_sqmuxa_1 (.A(un1_sersta65), .B(
        ack_1_sqmuxa_1_net_1), .C(pedetect_net_1), .D(
        \sercon[6]_net_1 ), .Y(serdat_1_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'h0013) )  \fsmmod_RNO[4]  (.A(\fsmmod[2]_net_1 ), 
        .B(\fsmmod_ns_i_0_0[4]_net_1 ), .C(N_213), .D(N_398), .Y(
        N_1013_i_0));
    CFG3 #( .INIT(8'h40) )  
        \SDAO_int_write_proc.un1_sersta65_1_2_1_a2_0  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[3]_net_1 ), .Y(N_1235));
    SLE \SCLI_ff_reg[2]  (.D(N_294_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[2]_net_1 ));
    CFG4 #( .INIT(16'hB0C0) )  \indelay_4[1]  (.A(\indelay[2]_net_1 ), 
        .B(\indelay[0]_net_1 ), .C(\fsmsync[3]_net_1 ), .D(
        \indelay[1]_net_1 ), .Y(\indelay_4[1]_net_1 ));
    CFG4 #( .INIT(16'h000D) )  \fsmsync_RNO[3]  (.A(N_973), .B(
        \fsmsync[3]_net_1 ), .C(\fsmsync_ns_i_0[3]_net_1 ), .D(N_990), 
        .Y(N_959_i_0));
    CFG4 #( .INIT(16'h0040) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_0  (.A(
        \fsmsta[4]_net_1 ), .B(fsmsta_9_0_372_i_0_a2_0_1), .C(
        fsmsta_9_0_372_i_0_a2_0_0), .D(N_356), .Y(N_441));
    CFG2 #( .INIT(4'h4) )  \fsmmod_ns_0_0_a2_0_2[5]  (.A(SDAInt_net_1), 
        .B(\fsmmod[0]_net_1 ), .Y(\fsmmod_ns_0_0_a2_0[5]_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  \sersta_write_proc.sersta_3_0[3]  (.A(
        N_289), .B(\sersta_3_0_1[3] ), .C(\fsmsta[3]_net_1 ), .D(N_549)
        , .Y(\sersta_3[3] ));
    SLE \fsmsync[3]  (.D(N_959_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  adrcomp_RNIH4RF (.A(counter_PRESETN_1), .B(
        adrcomp_net_1), .Y(fsmsta_m2_e_0));
    SLE \PCLK_count2[1]  (.D(\PCLK_count2_4[1]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\PCLK_count2[1]_net_1 ));
    CFG4 #( .INIT(16'hFFEA) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_i  (
        .A(fsmsta_9_2_342_i_i_0), .B(fsmsta_m2_e_0), .C(N_117), .D(
        N_449), .Y(N_94));
    CFG4 #( .INIT(16'h078F) )  
        \fsmsta_sync_proc.fsmsta_9_0_o2_1_2_1[0]  (.A(pedetect_net_1), 
        .B(framesync24), .C(N_543), .D(\fsmsta_9_0_a2_4_0[0] ), .Y(
        \fsmsta_9_0_o2_1_2_1[0] ));
    CFG4 #( .INIT(16'h0E04) )  \sersta_write_proc.sersta_3_0_1[1]  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(N_361), .D(N_393)
        , .Y(\sersta_3_0_1[1] ));
    CFG4 #( .INIT(16'h0040) )  \serdat_write_proc.un4_PRDATA  (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(controlReg14_3), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .D(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(un4_PRDATA));
    CFG4 #( .INIT(16'h1110) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_1  (.A(pedetect_net_1), 
        .B(counter_PRESETN_1), .C(N_509), .D(fsmsta_9_0_372_i_0_o2_1_4)
        , .Y(N_442));
    CFG4 #( .INIT(16'hFFF4) )  \fsmsta_sync_proc.fsmsta_9_0[4]  (.A(
        N_356), .B(\fsmsta_9_0_a2_1_2[4] ), .C(\fsmsta_9_0_3[4] ), .D(
        \fsmsta_9_0_1[4] ), .Y(\fsmsta_9[4] ));
    CFG4 #( .INIT(16'h1230) )  \PCLK_count2_4[1]  (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN_net_1), .C(
        \PCLK_count2[1]_net_1 ), .D(\PCLK_count2[0]_net_1 ), .Y(
        \PCLK_count2_4[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[3]  (.A(
        serdat4), .B(serdat_2), .C(CoreAPB3_0_APBmslave0_PWDATA[3]), 
        .Y(\serdat_19[3] ));
    CFG3 #( .INIT(8'hF4) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1_5[2]  (
        .A(N_355), .B(N_255), .C(\fsmsta_9_0_o2_1_2[2] ), .Y(
        \fsmsta_9_0_o2_1_4[2] ));
    CFG2 #( .INIT(4'hE) )  \PCLK_counter1_proc.PCLK_count1_4_i_o2[1]  
        (.A(counter_PRESETN_net_1), .B(\PCLK_count1[3]_net_1 ), .Y(
        N_238));
    CFG3 #( .INIT(8'hEF) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_3  
        (.A(\fsmmod[0]_net_1 ), .B(\fsmmod[5]_net_1 ), .C(
        un1_framesync24), .Y(N_419));
    CFG4 #( .INIT(16'hFFF2) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_1_1  (.A(
        fsmsta_9_0_372_i_0_a2_12_0), .B(N_364), .C(N_504), .D(N_507), 
        .Y(fsmsta_9_0_372_i_0_o2_1_1));
    CFG4 #( .INIT(16'h0008) )  \fsmmod_ns_0_0_a2_0[1]  (.A(
        SDAInt_net_1), .B(\fsmmod[0]_net_1 ), .C(N_398), .D(N_200), .Y(
        N_297));
    SLE busfree (.D(\fsmdet_i_0[3] ), .CLK(GL0_INST), .EN(un1_fsmdet), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(busfree_net_1));
    CFG4 #( .INIT(16'hDCCC) )  \fsmmod_ns_0_0[3]  (.A(N_398), .B(N_298)
        , .C(\fsmmod[3]_net_1 ), .D(N_407), .Y(\fsmmod_ns[3] ));
    SLE \PCLK_count1[2]  (.D(N_342_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[2]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \fsmsta_sync_proc.fsmsta_9_0_m2_1[4]  (.A(
        ack_net_1), .B(\fsmsta[4]_net_1 ), .C(N_129), .Y(N_410));
    CFG4 #( .INIT(16'h0800) )  \fsmmod_ns_0_0_a2[3]  (.A(
        \fsmmod_ns_0_0_a2_1[3] ), .B(N_162), .C(N_185), .D(
        un1_framesync_2), .Y(N_298));
    CFG4 #( .INIT(16'h0010) )  \PRDATA_0_iv_0_RNO_0[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(\sercon[4]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(sercon_m2_e_0_1));
    CFG4 #( .INIT(16'hCCCD) )  \fsmsync_ns_i_1[6]  (.A(un1_framesync_2)
        , .B(\fsmsync_ns_i_0[6]_net_1 ), .C(\fsmsync[6]_net_1 ), .D(
        \fsmsync[5]_net_1 ), .Y(\fsmsync_ns_i_1[6]_net_1 ));
    SLE \sercon[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[6]_net_1 ));
    SLE SDAO_int (.D(N_1272), .CLK(GL0_INST), .EN(
        SDAO_int_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\COREI2C_0_0_SDAO[0] ));
    CFG3 #( .INIT(8'hFE) )  
        \PCLK_counter1_proc.PCLK_count17_1.CO3_i_o2  (.A(
        \PCLK_count1[1]_net_1 ), .B(\PCLK_count1[0]_net_1 ), .C(
        \PCLK_count1[2]_net_1 ), .Y(N_220));
    CFG4 #( .INIT(16'h82D7) )  \sersta_write_proc.sersta_3_0_m2[2]  (
        .A(N_361), .B(N_358), .C(\fsmsta[2]_net_1 ), .D(N_393), .Y(
        N_414));
    CFG3 #( .INIT(8'hF8) )  \SDAO_int_write_proc.SDAO_int_6_0_312  (.A(
        SDAO_int_6_0_312_a5_0), .B(N_1289), .C(SDAO_int_6_0_312_1), .Y(
        N_1272));
    CFG2 #( .INIT(4'h4) )  \fsmsync_sync_proc.un1_sersta69_1_a5_0_0  (
        .A(\fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_492));
    CFG3 #( .INIT(8'hE0) )  \fsmmod_ns_i_0_a2_0_2[2]  (.A(N_364), .B(
        N_355), .C(un1_framesync_2), .Y(
        \fsmmod_ns_i_0_a2_0_2[2]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_2  
        (.A(\fsmmod[6]_net_1 ), .B(\fsmmod[1]_net_1 ), .C(
        \fsmdet[3]_net_1 ), .Y(N_443));
    CFG2 #( .INIT(4'h7) )  \fsmsta_sync_proc.fsmsta_9_0_o2_5[4]  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_358));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[2]  (.A(
        serdat4), .B(\serdat[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .Y(\serdat_19[2] ));
    CFG2 #( .INIT(4'h4) )  nedetect_0_sqmuxa_0_a2 (.A(N_262), .B(
        SCLInt_net_1), .Y(nedetect_0_sqmuxa));
    CFG4 #( .INIT(16'hB333) )  \fsmsta_sync_proc.fsmsta_9_0_0[4]  (.A(
        N_129), .B(N_221), .C(framesync24), .D(\fsmsta_9_0_a2_2_2[4] ), 
        .Y(\fsmsta_9_0_0[4] ));
    CFG4 #( .INIT(16'h0307) )  \fsmmod_ns_i_0_a2[2]  (.A(
        \fsmmod[1]_net_1 ), .B(nedetect_net_1), .C(\fsmmod[2]_net_1 ), 
        .D(\fsmmod[6]_net_1 ), .Y(N_452));
    CFG4 #( .INIT(16'hF1F0) )  \fsmsta_sync_proc.fsmsta_9_0_o2_3[0]  (
        .A(\fsmsta[2]_net_1 ), .B(ack_net_1), .C(
        \fsmsta_9_0_o2_3_0[0] ), .D(N_542), .Y(N_400));
    CFG4 #( .INIT(16'hEA00) )  \fsmdet_RNO[6]  (.A(\fsmdet[5]_net_1 ), 
        .B(\fsmdet[6]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_881_i_0));
    CFG2 #( .INIT(4'h1) )  \sercon_write_proc.sercon_9_0_0_a0_0[3]  (
        .A(CoreAPB3_0_APBmslave0_PADDR[8]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(un12_PSELi_0));
    CFG4 #( .INIT(16'h5410) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_4  
        (.A(counter_PRESETN_1), .B(framesync24), .C(N_554), .D(N_551), 
        .Y(fsmsta_9_0_372_i_0_4));
    CFG3 #( .INIT(8'hFB) )  \sercon_write_proc.sercon_9_i_o2[4]  (.A(
        N_372), .B(\sercon[4]_net_1 ), .C(N_527), .Y(N_418));
    CFG3 #( .INIT(8'h10) )  \PRDATA_0_iv_0_RNO[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(sercon_m2_e_1), .Y(
        \sercon_m[3] ));
    SLE \serdat[1]  (.D(\serdat_19[1] ), .CLK(GL0_INST), .EN(
        un1_N_9_mux_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\serdat[1]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \sercon_RNIIC4A2[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(sercon_m2_e_3_1), .Y(
        \sercon_m[1] ));
    CFG3 #( .INIT(8'h08) )  SDAO_int_1_sqmuxa_3 (.A(N_359), .B(
        SDAO_int_1_sqmuxa_1_net_1), .C(\fsmmod[1]_net_1 ), .Y(
        SDAO_int_1_sqmuxa_3_net_1));
    CFG4 #( .INIT(16'hFCDD) )  \fsmsta_sync_proc.fsmsta_9_0_o2_2[4]  (
        .A(N_361), .B(N_527), .C(N_410), .D(framesync24), .Y(N_228));
    CFG2 #( .INIT(4'hE) )  
        \SDAO_int_write_proc.un1_sersta65_1_2_0_o2_0  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[1]_net_1 ), .Y(N_364));
    CFG4 #( .INIT(16'h4EE4) )  
        \framesync_write_proc.framesync_6_enl[0]  (.A(framesync_6_e2), 
        .B(\framesync_6_m2[3] ), .C(\framesync[0]_net_1 ), .D(
        un1_nedetect), .Y(\framesync_6[0] ));
    CFG2 #( .INIT(4'h7) )  \SCLInt_write_proc.un1_SCLInt5_0  (.A(N_262)
        , .B(pedetect_0_sqmuxa_3), .Y(un1_SCLInt5));
    CFG3 #( .INIT(8'h08) )  un14_counter_PRESETN (.A(
        \COREI2C_0_0_SCLO[0] ), .B(\fsmmod[4]_net_1 ), .C(SCLInt_net_1)
        , .Y(un14_counter_PRESETN_net_1));
    CFG4 #( .INIT(16'hFFAE) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_o2_12_1  (.A(ack_net_1), 
        .B(un1_ack_1_0), .C(N_244), .D(N_527), .Y(
        fsmsta_9_0_372_i_0_o2_12_1));
    CFG4 #( .INIT(16'hF2F0) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0_3  
        (.A(counter_PRESETN_1), .B(adrcomp_net_1), .C(
        fsmsta_9_0_372_i_0_2), .D(N_419), .Y(fsmsta_9_0_372_i_0_3));
    CFG2 #( .INIT(4'h2) )  \fsmmod_ns_0_0_a2_0_0[5]  (.A(
        \fsmmod[5]_net_1 ), .B(sclscl_net_1), .Y(
        \fsmmod_ns_0_0_a2_0_0[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \sersta_write_proc.sersta_3_0_a2_1[4]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(sersta77_2));
    CFG4 #( .INIT(16'h0008) )  \fsmsta_sync_proc.fsmsta_9_0_a2_16[0]  
        (.A(SDAInt_net_1), .B(\fsmsta[1]_net_1 ), .C(\fsmsta[2]_net_1 )
        , .D(N_355), .Y(N_497));
    CFG3 #( .INIT(8'h40) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_13  (.A(N_355), .B(
        framesync24), .C(N_140_i), .Y(N_499));
    CFG4 #( .INIT(16'h0E00) )  \fsmdet_RNO[3]  (.A(\fsmdet[1]_net_1 ), 
        .B(\fsmdet[6]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_875_i_0));
    CFG3 #( .INIT(8'h02) )  \fsmsync_RNO[1]  (.A(\fsmsync[0]_net_1 ), 
        .B(SCLInt_net_1), .C(N_985), .Y(N_955_i_0));
    CFG4 #( .INIT(16'h8001) )  \SDAInt_write_proc.un1_SDAInt5_0  (.A(
        \SDAI_ff_reg[3]_net_1 ), .B(\SDAI_ff_reg[2]_net_1 ), .C(
        \SDAI_ff_reg[1]_net_1 ), .D(\SDAI_ff_reg[0]_net_1 ), .Y(
        un1_SDAInt5));
    CFG3 #( .INIT(8'h82) )  \indelay_4[0]  (.A(\fsmsync[3]_net_1 ), .B(
        fsmsync_nxt35), .C(\indelay[0]_net_1 ), .Y(
        \indelay_4[0]_net_1 ));
    CFG3 #( .INIT(8'hF7) )  \fsmsta_sync_proc.fsmsta_9_0_o2_6[4]  (.A(
        \fsmsta[2]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(SDAInt_net_1)
        , .Y(N_401));
    SLE \fsmsync[5]  (.D(N_963_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[5]_net_1 ));
    CFG3 #( .INIT(8'h75) )  \fsmsync_ns_i_o3[2]  (.A(
        \fsmsync[2]_net_1 ), .B(PCLKint_ff_net_1), .C(PCLKint_net_1), 
        .Y(N_979));
    CFG3 #( .INIT(8'hE4) )  \serdat_write_proc.serdat_19[4]  (.A(
        serdat4), .B(\serdat[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .Y(\serdat_19[4] ));
    CFG4 #( .INIT(16'hFFFB) )  \fsmsta_sync_proc.fsmsta_9_0_o2_1[0]  (
        .A(N_490), .B(\fsmsta_9_0_o2_1_2_1[0] ), .C(N_400), .D(
        \fsmsta_9_0_o2_1_1[0] ), .Y(N_353));
    CFG4 #( .INIT(16'hA800) )  \fsmsta_sync_proc.fsmsta_9_0_a2_1_2[4]  
        (.A(\fsmsta_9_0_a2_2_0[4] ), .B(N_374), .C(
        \COREI2C_0_0_SDAO[0] ), .D(N_129), .Y(\fsmsta_9_0_a2_1_2[4] ));
    CFG3 #( .INIT(8'hAB) )  \sercon_write_proc.sercon_9_0_o2[3]  (.A(
        adrcomp_net_1), .B(\fsmmod[5]_net_1 ), .C(\fsmmod[0]_net_1 ), 
        .Y(N_370));
    CFG4 #( .INIT(16'hF8FA) )  \fsmsync_ns_0_1[0]  (.A(SCLInt_net_1), 
        .B(\fsmsync[4]_net_1 ), .C(N_985), .D(N_980), .Y(
        \fsmsync_ns_0_1[0]_net_1 ));
    CFG4 #( .INIT(16'hCCAC) )  ack_RNO (.A(ack_10_u_yy), .B(
        ack_10_u_xx), .C(un1_serdat_2_sqmuxa_1_tz), .D(serdat4), .Y(
        ack_10));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_RNO[2]  (.A(\sercon[6]_net_1 ), 
        .B(\SDAI_ff_reg[1]_net_1 ), .Y(N_66_i_0));
    CFG2 #( .INIT(4'hE) )  
        \fsmsync_sync_proc.un1_sersta69_1_a5_2_2_0_o2  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .Y(N_394));
    CFG3 #( .INIT(8'h04) )  \sercon_write_proc.un1_PRDATA  (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(un1_WEn_0), .C(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(un1_PRDATA));
    CFG4 #( .INIT(16'hCC80) )  \fsmsync_ns_0_o3_0_a2[0]  (.A(
        \fsmmod[1]_net_1 ), .B(N_438_1), .C(\fsmmod[2]_net_1 ), .D(
        \fsmmod[3]_net_1 ), .Y(N_438));
    CFG3 #( .INIT(8'hD8) )  \SDAO_int_write_proc.un1_sersta58_0_m2  (
        .A(\fsmsta[2]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \fsmsta[4]_net_1 ), .Y(N_365));
    CFG4 #( .INIT(16'hFFFE) )  \fsmsync_sync_proc.un1_sersta69_1  (.A(
        N_1235), .B(sersta77_2), .C(N_1236), .D(N_466), .Y(
        un1_sersta69));
    CFG3 #( .INIT(8'h20) )  un14_PRDATA_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(un14_PRDATA_0_net_1));
    SLE \sersta[2]  (.D(\sersta_3[2] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[2]_net_1 ));
    CFG4 #( .INIT(16'h0220) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_0_a2_23  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \COREI2C_0_0_SDAO[0] ), .D(\fsmsta[0]_net_1 ), .Y(N_504));
    CFG4 #( .INIT(16'hFBF3) )  \sersta_write_proc.sersta_3_0[1]  (.A(
        N_374), .B(COREI2C_0_0_INT[0]), .C(\sersta_3_0_1[1] ), .D(
        N_361), .Y(\sersta_3[1] ));
    CFG4 #( .INIT(16'h0010) )  ack_1_sqmuxa_1 (.A(\fsmdet[3]_net_1 ), 
        .B(COREI2C_0_0_INT[0]), .C(un1_sersta65_1), .D(un1_sersta58_0), 
        .Y(ack_1_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'hE0A0) )  \indelay_4[2]  (.A(\indelay[2]_net_1 ), 
        .B(\indelay[0]_net_1 ), .C(\fsmsync[3]_net_1 ), .D(
        \indelay[1]_net_1 ), .Y(\indelay_4[2]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \fsmsta_sync_proc.fsmsta_9_0_o2_3_0[2]  (.A(
        SDAInt_net_1), .B(sercon_2), .Y(\fsmsta_9_0_o2_3_0[2] ));
    CFG2 #( .INIT(4'h8) )  \sersta_write_proc.sersta_3_0_a2[2]  (.A(
        N_524), .B(\fsmsta[1]_net_1 ), .Y(N_543));
    CFG4 #( .INIT(16'h2000) )  
        \serdat_write_proc.un4_PRDATA_1_RNIJ9E51  (.A(
        \serdat[1]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[0]), .C(
        un4_PRDATA_1), .D(controlReg14_3), .Y(\serdat_m[1] ));
    
endmodule


module COREI2C_Z3(
       COREI2C_0_0_SDAO_i,
       COREI2C_0_0_SCLO_i,
       COREI2C_0_0_INT,
       CoreAPB3_0_APBmslave0_PADDR,
       CoreAPB3_0_APBmslave0_PRDATA_m_1,
       CoreAPB3_0_APBmslave0_PRDATA_m_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_2,
       TRIG_c,
       gpin3_m_2_0,
       GPOUT_reg,
       gpin3_m,
       CoreAPB3_0_APBmslave1_PRDATA_m,
       CoreAPB3_0_APBmslave0_PWDATA,
       sercon_0,
       sercon_2,
       serdat_2,
       serdat_0,
       CoreAPB3_0_APBmslave0_PRDATA_m_0_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_4,
       CoreAPB3_0_APBmslave0_PRDATA_m_2_d0,
       CoreAPB3_0_APBmslave0_PRDATA_m_3,
       CoreAPB3_0_APBmslave0_PRDATA_m_5,
       un12_PSELi,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       r_N_4_mux,
       N_97_1,
       controlReg14_3,
       un4_PRDATA_1,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       un1_WEn_1,
       BIBUF_COREI2C_0_0_SCL_IO_Y,
       BIBUF_COREI2C_0_0_SDA_IO_Y,
       un1_WEn_0,
       un14_PRDATA,
       un1_PRDATA,
       un4_PRDATA,
       CoreAPB3_0_APBmslave0_PSELx,
       GPOUT_reg40_2,
       CoreAPB3_0_APBmslave1_PSELx,
       GPOUT_reg40
    );
output [0:0] COREI2C_0_0_SDAO_i;
output [0:0] COREI2C_0_0_SCLO_i;
output [0:0] COREI2C_0_0_INT;
input  [8:0] CoreAPB3_0_APBmslave0_PADDR;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_1;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_0;
output [7:7] CoreAPB3_0_APBmslave0_PRDATA_m_2;
input  [0:0] TRIG_c;
input  [1:1] gpin3_m_2_0;
input  [1:1] GPOUT_reg;
input  [1:1] gpin3_m;
output [1:0] CoreAPB3_0_APBmslave1_PRDATA_m;
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output sercon_0;
output sercon_2;
output serdat_2;
output serdat_0;
output CoreAPB3_0_APBmslave0_PRDATA_m_0_d0;
output CoreAPB3_0_APBmslave0_PRDATA_m_4;
output CoreAPB3_0_APBmslave0_PRDATA_m_2_d0;
output CoreAPB3_0_APBmslave0_PRDATA_m_3;
output CoreAPB3_0_APBmslave0_PRDATA_m_5;
output un12_PSELi;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  r_N_4_mux;
output N_97_1;
output controlReg14_3;
output un4_PRDATA_1;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
output un1_WEn_1;
input  BIBUF_COREI2C_0_0_SCL_IO_Y;
input  BIBUF_COREI2C_0_0_SDA_IO_Y;
output un1_WEn_0;
output un14_PRDATA;
output un1_PRDATA;
output un4_PRDATA;
input  CoreAPB3_0_APBmslave0_PSELx;
input  GPOUT_reg40_2;
input  CoreAPB3_0_APBmslave1_PSELx;
input  GPOUT_reg40;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    COREI2CREAL_Z4 \I2C_NUM_GENERATION[0].ui2c  (.COREI2C_0_0_SDAO_i({
        COREI2C_0_0_SDAO_i[0]}), .COREI2C_0_0_SCLO_i({
        COREI2C_0_0_SCLO_i[0]}), .COREI2C_0_0_INT({COREI2C_0_0_INT[0]})
        , .CoreAPB3_0_APBmslave0_PADDR({CoreAPB3_0_APBmslave0_PADDR[8], 
        CoreAPB3_0_APBmslave0_PADDR[7], CoreAPB3_0_APBmslave0_PADDR[6], 
        CoreAPB3_0_APBmslave0_PADDR[5], CoreAPB3_0_APBmslave0_PADDR[4], 
        CoreAPB3_0_APBmslave0_PADDR[3], CoreAPB3_0_APBmslave0_PADDR[2], 
        CoreAPB3_0_APBmslave0_PADDR[1], CoreAPB3_0_APBmslave0_PADDR[0]})
        , .CoreAPB3_0_APBmslave0_PRDATA_m_1({
        CoreAPB3_0_APBmslave0_PRDATA_m_1[7]}), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_0({
        CoreAPB3_0_APBmslave0_PRDATA_m_0[7]}), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2({
        CoreAPB3_0_APBmslave0_PRDATA_m_2[7]}), .TRIG_c({TRIG_c[0]}), 
        .gpin3_m_2_0({gpin3_m_2_0[1]}), .GPOUT_reg({GPOUT_reg[1]}), 
        .gpin3_m({gpin3_m[1]}), .CoreAPB3_0_APBmslave1_PRDATA_m({
        CoreAPB3_0_APBmslave1_PRDATA_m[1], 
        CoreAPB3_0_APBmslave1_PRDATA_m[0]}), 
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .sercon_0(sercon_0), 
        .sercon_2(sercon_2), .serdat_2(serdat_2), .serdat_0(serdat_0), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_0_d0(
        CoreAPB3_0_APBmslave0_PRDATA_m_0_d0), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_4(
        CoreAPB3_0_APBmslave0_PRDATA_m_4), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2_d0(
        CoreAPB3_0_APBmslave0_PRDATA_m_2_d0), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_3(
        CoreAPB3_0_APBmslave0_PRDATA_m_3), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_5(
        CoreAPB3_0_APBmslave0_PRDATA_m_5), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .r_N_4_mux(
        r_N_4_mux), .N_97_1(N_97_1), .controlReg14_3(controlReg14_3), 
        .un4_PRDATA_1(un4_PRDATA_1), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .un1_WEn_1(un1_WEn_1), 
        .BIBUF_COREI2C_0_0_SCL_IO_Y(BIBUF_COREI2C_0_0_SCL_IO_Y), 
        .BIBUF_COREI2C_0_0_SDA_IO_Y(BIBUF_COREI2C_0_0_SDA_IO_Y), 
        .un1_WEn_0(un1_WEn_0), .un14_PRDATA(un14_PRDATA), .un1_PRDATA(
        un1_PRDATA), .un4_PRDATA(un4_PRDATA), 
        .CoreAPB3_0_APBmslave0_PSELx(CoreAPB3_0_APBmslave0_PSELx), 
        .un12_PSELi(un12_PSELi), .GPOUT_reg40_2(GPOUT_reg40_2), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .GPOUT_reg40(GPOUT_reg40));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0001) )  \I2C_NUM_PSELi_GEN[0].un12_PSELi  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[8]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(un12_PSELi));
    
endmodule


module CoreResetP_Z7(
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       SYSRESET_POR,
       mss_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N
    );
output MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  SYSRESET_POR;
input  mss_sb_MSS_TMP_0_MSS_RESET_N_M2F;
input  mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N;

    wire MSS_HPMS_READY_int_net_1, mss_ready_select_net_1, VCC_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        GND_net_1, mss_ready_state_net_1, RESET_N_M2F_clk_base_net_1, 
        POWER_ON_RESET_N_q1_net_1, RESET_N_M2F_q1_net_1, 
        FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, MSS_HPMS_READY_int_4_net_1;
    
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(RESET_N_M2F_clk_base_net_1));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_clk_base_net_1));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        mss_ready_select4_net_1), .ALn(POWER_ON_RESET_N_clk_base_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(mss_ready_select_net_1));
    CLKINT MSS_HPMS_READY_int_RNI5CTC_inst_1 (.A(
        MSS_HPMS_READY_int_net_1), .Y(MSS_HPMS_READY_int_RNI5CTC));
    GND GND (.Y(GND_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        RESET_N_M2F_clk_base_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_q1_net_1));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_q1_net_1));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Rx_async_1s_0s_1s_2s(
       rx_byte,
       rx_state,
       controlReg2,
       clear_parity_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       BT_TX_c,
       CoreUARTapb_2_0_PARITY_ERR,
       stop_strobe,
       CoreUARTapb_2_0_FRAMING_ERR,
       clear_parity_en,
       fifo_write
    );
output [7:0] rx_byte;
output [1:0] rx_state;
input  [2:0] controlReg2;
input  clear_parity_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  baud_clock;
input  BT_TX_c;
output CoreUARTapb_2_0_PARITY_ERR;
output stop_strobe;
output CoreUARTapb_2_0_FRAMING_ERR;
output clear_parity_en;
output fifo_write;

    wire clear_parity_reg_i_0, \rx_bit_cnt[0]_net_1 , VCC_net_1, 
        \rx_bit_cnt_4[0] , GND_net_1, \rx_bit_cnt[1]_net_1 , 
        \rx_bit_cnt_4[1] , \rx_bit_cnt[2]_net_1 , \rx_bit_cnt_4[2] , 
        \rx_bit_cnt[3]_net_1 , \rx_bit_cnt_4[3] , \samples[1]_net_1 , 
        \samples[2]_net_1 , \rx_shift[0]_net_1 , \rx_shift_11[0] , 
        un1_samples7_1_0_net_1, \rx_shift[1]_net_1 , \rx_shift_11[1] , 
        \rx_shift[2]_net_1 , \rx_shift_11[2] , \rx_shift[3]_net_1 , 
        \rx_shift_11[3] , \rx_shift[4]_net_1 , \rx_shift_11[4] , 
        \rx_shift[5]_net_1 , \rx_shift_11[5] , \rx_shift[6]_net_1 , 
        \rx_shift_11[6] , \rx_shift[7]_net_1 , \rx_shift_11[7] , 
        \rx_shift[8]_net_1 , \rx_shift_11[8] , 
        \receive_count[0]_net_1 , \receive_count_3[0] , 
        \receive_count[1]_net_1 , \receive_count_3[1] , 
        \receive_count[2]_net_1 , \receive_count_3[2] , 
        \receive_count[3]_net_1 , \receive_count_3[3] , 
        clear_parity_en_9, \rx_byte_2[7] , \samples[0]_net_1 , N_310, 
        parity_err_1_sqmuxa_i_0, rx_parity_calc_net_1, 
        rx_parity_calc_4, framing_error_int_net_1, 
        framing_error_int_0_sqmuxa_net_1, framing_error_int_2_sqmuxa, 
        framing_error_1_sqmuxa_i_0, N_233_i_0, \rx_state_ns[0] , 
        clear_parity_en_9_i_0, N_238_3, rx_state19_li, CO1, 
        rx_bit_cnt_0_sqmuxa, un1_parity_err_0_sqmuxa_2_1_1_net_1, 
        un1_parity_err_0_sqmuxa_2_1_net_1, un1_parity_err31_0_net_1, 
        N_238_1, N_242, framing_error_int_0_sqmuxa_1_net_1, rx_state10, 
        rx_state19_0, framing_error_int5, rx_state19_NE_1, 
        rx_bit_cnt_1_sqmuxa, rx_parity_calc4, \rx_shift_9[8] , 
        \rx_shift_9[7] , \rx_shift_9[6] , receive_count8;
    
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_samples7_1_0 (.A(baud_clock), .B(
        N_238_3), .C(rx_bit_cnt_0_sqmuxa), .Y(un1_samples7_1_0_net_1));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[0]));
    CFG4 #( .INIT(16'h8000) )  framing_error_int_0_sqmuxa (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        framing_error_int5), .D(framing_error_int_0_sqmuxa_1_net_1), 
        .Y(framing_error_int_0_sqmuxa_net_1));
    SLE \receive_count[1]  (.D(\receive_count_3[1] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[1]_net_1 ));
    SLE \rx_shift[7]  (.D(\rx_shift_11[7] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \rx_par_calc.rx_parity_calc4  (.A(N_238_3), 
        .B(controlReg2[1]), .Y(rx_parity_calc4));
    CFG4 #( .INIT(16'h1441) )  
        \make_parity_err.parity_err_12_iv_0_111_a2  (.A(
        clear_parity_reg), .B(framing_error_int5), .C(
        rx_parity_calc_net_1), .D(controlReg2[2]), .Y(N_310));
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[0]_net_1 ));
    CFG4 #( .INIT(16'h72F0) )  \receive_shift.rx_shift_11_RNO[8]  (.A(
        controlReg2[1]), .B(framing_error_int5), .C(
        \rx_shift[8]_net_1 ), .D(controlReg2[0]), .Y(\rx_shift_9[8] ));
    CFG3 #( .INIT(8'h40) )  
        \receive_full_indicator.clear_parity_en_9_0_a3  (.A(
        rx_state19_li), .B(rx_state[0]), .C(baud_clock), .Y(
        clear_parity_en_9));
    CFG2 #( .INIT(4'h1) )  \rcv_cnt.receive_count_3[0]  (.A(
        receive_count8), .B(\receive_count[0]_net_1 ), .Y(
        \receive_count_3[0] ));
    CFG1 #( .INIT(2'h1) )  framing_error_RNO (.A(clear_parity_reg), .Y(
        clear_parity_reg_i_0));
    CFG3 #( .INIT(8'h06) )  \rcv_cnt.receive_count_3[1]  (.A(
        \receive_count[1]_net_1 ), .B(\receive_count[0]_net_1 ), .C(
        receive_count8), .Y(\receive_count_3[1] ));
    CFG3 #( .INIT(8'h14) )  \rcv_cnt.receive_count_3[2]  (.A(
        receive_count8), .B(\receive_count[2]_net_1 ), .C(N_238_1), .Y(
        \receive_count_3[2] ));
    CFG3 #( .INIT(8'h04) )  rx_bit_cnt_0_sqmuxa_0_a3 (.A(rx_state[1]), 
        .B(baud_clock), .C(rx_state[0]), .Y(rx_bit_cnt_0_sqmuxa));
    CFG4 #( .INIT(16'h90F6) )  \receive_shift.rx_shift_9_u[7]  (.A(
        controlReg2[0]), .B(controlReg2[1]), .C(N_242), .D(
        framing_error_int5), .Y(\rx_shift_9[7] ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[0]  (.A(
        \rx_shift[1]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(\receive_count_3[3] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[4]));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[8]  (.A(
        rx_state[1]), .B(\rx_shift_9[8] ), .C(rx_state[0]), .Y(
        \rx_shift_11[8] ));
    SLE rx_parity_calc (.D(rx_parity_calc_4), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_parity_calc_net_1));
    SLE \rx_bit_cnt[2]  (.D(\rx_bit_cnt_4[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[2]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[3]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(CO1), .D(
        rx_bit_cnt_0_sqmuxa), .Y(\rx_bit_cnt_4[3] ));
    CFG4 #( .INIT(16'h0002) )  \rcv_cnt.rx_state10_0_a3  (.A(
        \receive_count[3]_net_1 ), .B(\receive_count[2]_net_1 ), .C(
        \receive_count[1]_net_1 ), .D(\receive_count[0]_net_1 ), .Y(
        rx_state10));
    SLE \rx_bit_cnt[1]  (.D(\rx_bit_cnt_4[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[1]_net_1 ));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[7]  (.A(
        rx_state[1]), .B(\rx_shift_9[7] ), .C(rx_state[0]), .Y(
        \rx_shift_11[7] ));
    CFG3 #( .INIT(8'hAC) )  \receive_shift.rx_shift_9_0[7]  (.A(
        \rx_shift[8]_net_1 ), .B(\rx_shift[7]_net_1 ), .C(
        controlReg2[1]), .Y(N_242));
    CFG4 #( .INIT(16'hFFBD) )  \rcv_sm.rx_state19_NE_1  (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(
        \rx_bit_cnt[1]_net_1 ), .D(rx_state19_0), .Y(rx_state19_NE_1));
    SLE stop_strobe_inst_1 (.D(framing_error_int_2_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG4 #( .INIT(16'h0C2E) )  \rx_state_RNO[1]  (.A(rx_state[0]), .B(
        rx_state[1]), .C(N_238_3), .D(rx_state19_li), .Y(N_233_i_0));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[1]));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[2]  (.A(
        \rx_shift[3]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(\receive_count_3[2] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[2]_net_1 ));
    SLE clear_parity_en_1 (.D(clear_parity_en_9), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_en));
    CFG4 #( .INIT(16'h0180) )  un1_parity_err_0_sqmuxa_2_1 (.A(
        controlReg2[0]), .B(un1_parity_err_0_sqmuxa_2_1_1_net_1), .C(
        \rx_bit_cnt[3]_net_1 ), .D(\rx_bit_cnt[1]_net_1 ), .Y(
        un1_parity_err_0_sqmuxa_2_1_net_1));
    CFG4 #( .INIT(16'h8000) )  \un1_rx_bit_cnt_1.CO1  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        baud_clock), .D(N_238_3), .Y(CO1));
    SLE \rx_state[1]  (.D(N_233_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_state[1]));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[6]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h8000) )  \rx_state_ns_i_a3_0_3[1]  (.A(
        \receive_count[3]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[0]_net_1 ), .Y(
        N_238_3));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[4]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[3]  (.A(
        \rx_shift[4]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(\rx_byte_2[7] ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[7]));
    CFG4 #( .INIT(16'hFCED) )  \rcv_sm.rx_state19_NE  (.A(
        controlReg2[1]), .B(rx_state19_NE_1), .C(\rx_bit_cnt[1]_net_1 )
        , .D(controlReg2[0]), .Y(rx_state19_li));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[2]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(CO1), .Y(
        \rx_bit_cnt_4[2] ));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[3]));
    CFG2 #( .INIT(4'h8) )  rx_bit_cnt_1_sqmuxa_0_a3 (.A(N_238_3), .B(
        baud_clock), .Y(rx_bit_cnt_1_sqmuxa));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[2]));
    CFG2 #( .INIT(4'h8) )  \rcv_sm.rx_byte_2[7]  (.A(controlReg2[0]), 
        .B(\rx_shift[7]_net_1 ), .Y(\rx_byte_2[7] ));
    SLE parity_err (.D(N_310), .CLK(GL0_INST), .EN(
        parity_err_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_0_PARITY_ERR));
    SLE \rx_shift[6]  (.D(\rx_shift_11[6] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[6]_net_1 ));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[1]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[4]  (.A(
        \rx_shift[5]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[3]_net_1 ));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[6]  (.A(
        rx_state[1]), .B(\rx_shift_9[6] ), .C(rx_state[0]), .Y(
        \rx_shift_11[6] ));
    SLE framing_error_int (.D(framing_error_int_0_sqmuxa_net_1), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(framing_error_int_net_1));
    CFG3 #( .INIT(8'h69) )  \rcv_sm.rx_state19_0  (.A(controlReg2[1]), 
        .B(\rx_bit_cnt[0]_net_1 ), .C(controlReg2[0]), .Y(rx_state19_0)
        );
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_state[0]));
    CFG4 #( .INIT(16'h1101) )  \rcv_cnt.receive_count8  (.A(
        rx_state[0]), .B(rx_state[1]), .C(framing_error_int5), .D(
        rx_state10), .Y(receive_count8));
    SLE \samples[2]  (.D(BT_TX_c), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    CFG4 #( .INIT(16'h060C) )  \rcv_cnt.receive_count_3[3]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        receive_count8), .D(N_238_1), .Y(\receive_count_3[3] ));
    SLE \receive_count[0]  (.D(\receive_count_3[0] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[5]));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[5]  (.A(
        \rx_shift[6]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[5] ));
    CFG3 #( .INIT(8'hBF) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_i  (.A(
        rx_state19_li), .B(rx_state[0]), .C(baud_clock), .Y(
        clear_parity_en_9_i_0));
    CFG2 #( .INIT(4'h8) )  \rx_state_ns_i_a3_0[1]  (.A(N_238_3), .B(
        rx_state[1]), .Y(framing_error_int_2_sqmuxa));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[0]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(
        rx_bit_cnt_1_sqmuxa), .Y(\rx_bit_cnt_4[0] ));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[5]_net_1 ));
    CFG4 #( .INIT(16'hBA10) )  \rx_state_ns_0[0]  (.A(rx_state[0]), .B(
        rx_state[1]), .C(rx_state10), .D(rx_state19_li), .Y(
        \rx_state_ns[0] ));
    CFG2 #( .INIT(4'h7) )  un1_parity_err31_0 (.A(baud_clock), .B(
        controlReg2[1]), .Y(un1_parity_err31_0_net_1));
    SLE \rx_bit_cnt[0]  (.D(\rx_bit_cnt_4[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[0]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  framing_error_1_sqmuxa_i (.A(
        framing_error_int_net_1), .B(clear_parity_reg), .C(baud_clock), 
        .Y(framing_error_1_sqmuxa_i_0));
    CFG3 #( .INIT(8'h17) )  un1_parity_err_0_sqmuxa_2_1_1 (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(
        \rx_bit_cnt[0]_net_1 ), .Y(un1_parity_err_0_sqmuxa_2_1_1_net_1)
        );
    SLE \rx_shift[8]  (.D(\rx_shift_11[8] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \rx_state_ns_i_a3_0_1[1]  (.A(
        \receive_count[0]_net_1 ), .B(\receive_count[1]_net_1 ), .Y(
        N_238_1));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[1]  (.A(
        \rx_shift[2]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[1] ));
    CFG3 #( .INIT(8'h40) )  framing_error_int_0_sqmuxa_1 (.A(
        \receive_count[0]_net_1 ), .B(rx_state[1]), .C(
        \receive_count[1]_net_1 ), .Y(
        framing_error_int_0_sqmuxa_1_net_1));
    CFG3 #( .INIT(8'h17) )  \rx_filtered.m3  (.A(\samples[1]_net_1 ), 
        .B(\samples[0]_net_1 ), .C(\samples[2]_net_1 ), .Y(
        framing_error_int5));
    SLE framing_error (.D(clear_parity_reg_i_0), .CLK(GL0_INST), .EN(
        framing_error_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_0_FRAMING_ERR));
    CFG4 #( .INIT(16'hF0B1) )  \receive_shift.rx_shift_11_RNO[6]  (.A(
        controlReg2[1]), .B(framing_error_int5), .C(
        \rx_shift[7]_net_1 ), .D(controlReg2[0]), .Y(\rx_shift_9[6] ));
    CFG4 #( .INIT(16'hAEAA) )  parity_err_1_sqmuxa_i (.A(
        clear_parity_reg), .B(N_238_3), .C(un1_parity_err31_0_net_1), 
        .D(un1_parity_err_0_sqmuxa_2_1_net_1), .Y(
        parity_err_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'h2122) )  \rx_par_calc.rx_parity_calc_4_u  (.A(
        rx_parity_calc_net_1), .B(rx_state[1]), .C(framing_error_int5), 
        .D(rx_parity_calc4), .Y(rx_parity_calc_4));
    SLE \rx_bit_cnt[3]  (.D(\rx_bit_cnt_4[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[1]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        rx_bit_cnt_1_sqmuxa), .D(rx_bit_cnt_0_sqmuxa), .Y(
        \rx_bit_cnt_4[1] ));
    
endmodule


module mss_sb_CoreUARTapb_2_0_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] tx_hold_reg;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), .C_WEN(
        INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), 
        .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_ctrl_128(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_2353_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, \counter[0]_net_1 , 
        VCC_net_1, un1_counter_cry_0_Y_0, GND_net_1, 
        \counter[1]_net_1 , un1_counter_cry_1_0_S, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S, \counter[6]_net_1 , un1_counter_s_6_S, 
        \data_out_0[2] , \data_out_0[3] , \data_out_0[4] , 
        \data_out_0[5] , \data_out_0[6] , \data_out_0[7] , 
        \data_out_0[0] , \data_out_0[1] , \wr_pointer[1]_net_1 , 
        \wr_pointer_s[1] , \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_129_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_130_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        empty_4_net_1, full_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_130_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_2_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[2]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S), .Y(), .FCO(
        un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[3]));
    CFG4 #( .INIT(16'h7FFF) )  full_4_RNIGLBA (.A(\counter[0]_net_1 ), 
        .B(full_4_net_1), .C(\counter[6]_net_1 ), .D(
        \counter[4]_net_1 ), .Y(fifo_full_tx_i_0));
    SLE \counter[6]  (.D(un1_counter_s_6_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_129 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_129_FCO));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_4_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[4]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_129_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[5]));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_130 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_130_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIHRB7 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[6]));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_3_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[3]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_tx), .C(fifo_write_tx), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_0), 
        .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[4]_net_1 ), 
        .Y(fifo_empty_tx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_2353_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_1_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_5_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[5]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_2353_i_0 (.A(fifo_write_tx), .Y(
        N_2353_i_0_net_1));
    mss_sb_CoreUARTapb_2_0_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg({
        tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], 
        tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]})
        , .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_tx(fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(\counter[6]_net_1 ), 
        .FCI(un1_counter_cry_5), .S(un1_counter_s_6_S), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_256x8(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_0_fifo_ctrl_128 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.tx_dout_reg({
        tx_dout_reg[7], tx_dout_reg[6], tx_dout_reg[5], tx_dout_reg[4], 
        tx_dout_reg[3], tx_dout_reg[2], tx_dout_reg[1], tx_dout_reg[0]})
        , .tx_hold_reg({tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], 
        tx_hold_reg[4], tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], 
        tx_hold_reg[0]}), .fifo_write_tx(fifo_write_tx), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       controlReg2,
       fifo_read_tx,
       fifo_read_tx_i_0,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       xmit_pulse,
       BT_RX_c,
       CoreUARTapb_2_0_TXRDY,
       fifo_full_tx_i_0,
       xmit_clock,
       baud_clock,
       fifo_empty_tx
    );
input  [7:0] tx_dout_reg;
input  [2:0] controlReg2;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  xmit_pulse;
output BT_RX_c;
output CoreUARTapb_2_0_TXRDY;
input  fifo_full_tx_i_0;
input  xmit_clock;
input  baud_clock;
input  fifo_empty_tx;

    wire \tx_byte[4]_net_1 , VCC_net_1, N_133_i_0, GND_net_1, 
        \tx_byte[5]_net_1 , \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_122_i_0, \xmit_bit_sel[2]_net_1 , 
        N_124_i_0, \xmit_bit_sel[3]_net_1 , N_126_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , \tx_byte[2]_net_1 , 
        \tx_byte[3]_net_1 , tx_parity_net_1, tx_parity_5, 
        un1_tx_parity_1_sqmuxa_0_net_1, tx_4_iv_i_0, N_144_i_0, 
        \xmit_state_ns_i_0[6] , \xmit_state[6]_net_1 , 
        \xmit_state_ns[6] , \xmit_state[0]_net_1 , 
        \xmit_state_ns[0]_net_1 , \xmit_state[1]_net_1 , 
        \xmit_state[2]_net_1 , \xmit_state_ns[2]_net_1 , 
        \xmit_state[3]_net_1 , N_112_i_0, \xmit_state[4]_net_1 , 
        \xmit_state_ns[4]_net_1 , \xmit_state[5]_net_1 , 
        \xmit_state_ns[5]_net_1 , N_174, tx_2_u_am_1_1, tx_2_u_am, 
        tx_2_u_bm_1_1, tx_2_u_bm, tx_2, N_128_i, N_129, tx_3_i_m, 
        N_172, N_154;
    
    SLE tx_parity (.D(tx_parity_5), .CLK(GL0_INST), .EN(
        un1_tx_parity_1_sqmuxa_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_parity_net_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_0_TXRDY));
    CFG4 #( .INIT(16'h2000) )  \xmit_state_ns_a3[5]  (.A(
        \xmit_state[3]_net_1 ), .B(controlReg2[1]), .C(xmit_pulse), .D(
        N_172), .Y(N_154));
    CFG2 #( .INIT(4'h6) )  \xmit_state_ns_i_x2[3]  (.A(controlReg2[0]), 
        .B(\xmit_bit_sel[0]_net_1 ), .Y(N_128_i));
    SLE \xmit_state[3]  (.D(N_112_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[3]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \xmit_cnt.xmit_bit_sel_3_i_o2[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        N_129));
    CFG4 #( .INIT(16'h0031) )  \xmit_sel.tx_4_iv_i  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(tx_2), 
        .D(tx_3_i_m), .Y(tx_4_iv_i_0));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[0]_net_1 ));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[4]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_state_RNI879Q1[1]  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(
        xmit_pulse), .D(\xmit_state[6]_net_1 ), .Y(N_144_i_0));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNI169 (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[0]_net_1 ), .B(\xmit_bit_sel[1]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_122_i_0));
    CFG4 #( .INIT(16'h8000) )  un1_tx_parity_1_sqmuxa_0_a2 (.A(
        \xmit_state[3]_net_1 ), .B(xmit_clock), .C(baud_clock), .D(
        controlReg2[1]), .Y(N_174));
    VCC VCC (.Y(VCC_net_1));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[5]_net_1 ));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[5]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(tx_2_u_bm_1_1), 
        .D(\xmit_bit_sel[1]_net_1 ), .Y(tx_2_u_bm));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(
        xmit_pulse), .Y(\xmit_state_ns[2]_net_1 ));
    CFG4 #( .INIT(16'hDC50) )  \xmit_state_ns[4]  (.A(xmit_pulse), .B(
        N_172), .C(\xmit_state[4]_net_1 ), .D(N_174), .Y(
        \xmit_state_ns[4]_net_1 ));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_126_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[3]_net_1 ));
    SLE \xmit_bit_sel[2]  (.D(N_124_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \xmit_sel.tx_2_u_ns  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(tx_2_u_bm), .C(tx_2_u_am), .Y(
        tx_2));
    SLE tx (.D(tx_4_iv_i_0), .CLK(GL0_INST), .EN(N_144_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BT_RX_c));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[3]_net_1 ));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[7]_net_1 ));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_bm_1_1));
    CFG2 #( .INIT(4'hE) )  un1_tx_parity_1_sqmuxa_0 (.A(N_174), .B(
        \xmit_state[5]_net_1 ), .Y(un1_tx_parity_1_sqmuxa_0_net_1));
    CFG4 #( .INIT(16'hF7A0) )  \xmit_state_RNO[3]  (.A(xmit_pulse), .B(
        N_172), .C(\xmit_state[2]_net_1 ), .D(\xmit_state[3]_net_1 ), 
        .Y(N_112_i_0));
    CFG3 #( .INIT(8'h06) )  \xmit_par_calc.tx_parity_5  (.A(tx_2), .B(
        tx_parity_net_1), .C(\xmit_state[5]_net_1 ), .Y(tx_parity_5));
    CFG4 #( .INIT(16'h0040) )  \xmit_state_ns_i_a2[3]  (.A(
        \xmit_bit_sel[3]_net_1 ), .B(\xmit_bit_sel[2]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(N_128_i), .Y(N_172));
    CFG3 #( .INIT(8'h82) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_state[3]_net_1 ), .B(N_129), .C(\xmit_bit_sel[2]_net_1 ), 
        .Y(N_124_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_am_1_1));
    CFG4 #( .INIT(16'hFDEC) )  \xmit_state_ns[5]  (.A(xmit_pulse), .B(
        N_154), .C(\xmit_state[4]_net_1 ), .D(\xmit_state[5]_net_1 ), 
        .Y(\xmit_state_ns[5]_net_1 ));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[6]_net_1 ));
    CFG3 #( .INIT(8'h82) )  \xmit_sel.tx_4_iv_i_RNO  (.A(
        \xmit_state[4]_net_1 ), .B(controlReg2[2]), .C(tx_parity_net_1)
        , .Y(tx_3_i_m));
    SLE \xmit_bit_sel[1]  (.D(N_122_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[1]_net_1 ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[1]_net_1 ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(GL0_INST), 
        .EN(xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[2]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(tx_2_u_am_1_1), 
        .D(\xmit_bit_sel[1]_net_1 ), .Y(tx_2_u_am));
    CFG2 #( .INIT(4'h4) )  fifo_read_en0_1_i_a3 (.A(fifo_empty_tx), .B(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[6] ));
    SLE fifo_read_en0 (.D(\xmit_state_ns_i_0[6] ), .CLK(GL0_INST), .EN(
        N_144_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns[0]  (.A(fifo_empty_tx), 
        .B(xmit_pulse), .C(\xmit_state[5]_net_1 ), .D(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[0]_net_1 ));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[1]_net_1 ));
    SLE \xmit_state[4]  (.D(\xmit_state_ns[4]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[4]_net_1 ));
    CFG4 #( .INIT(16'h82A0) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_state[3]_net_1 ), .B(N_129), .C(\xmit_bit_sel[3]_net_1 ), 
        .D(\xmit_bit_sel[2]_net_1 ), .Y(N_126_i_0));
    CFG2 #( .INIT(4'h8) )  \xmit_state_RNIFJ9T[2]  (.A(xmit_pulse), .B(
        \xmit_state[2]_net_1 ), .Y(N_133_i_0));
    SLE \xmit_state[6]  (.D(\xmit_state_ns[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[6]_net_1 ));
    CFG2 #( .INIT(4'hB) )  fifo_read_en0_1_i_a3_i (.A(fifo_empty_tx), 
        .B(\xmit_state[0]_net_1 ), .Y(\xmit_state_ns_i_0[6] ));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Clock_gen_0s(
       controlReg1,
       controlReg2,
       xmit_clock,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       xmit_pulse
    );
input  [7:0] controlReg1;
input  [7:3] controlReg2;
output xmit_clock;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output baud_clock;
output xmit_pulse;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNIQ6LQ_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI89KCK[11]  (.A(
        VCC_net_1), .B(controlReg2[6]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[11] ), .FCI(\baud_cntr_cry[10] ), .S(
        \baud_cntr_s[11] ), .Y(), .FCO(\baud_cntr_cry[11] ));
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIRMIG2[0]  (.A(
        VCC_net_1), .B(controlReg1[0]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[0] ), .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), 
        .Y(), .FCO(\baud_cntr_cry[0] ));
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[1] ));
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[3] ));
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[3]_net_1 ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[9] ));
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNIQ6LQ_Y), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(baud_clock));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIQ03AE[7]  (.A(
        VCC_net_1), .B(controlReg1[7]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[7] ), .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] )
        , .Y(), .FCO(\baud_cntr_cry[7] ));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[7] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[5] ));
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIAJBI7[3]  (.A(
        VCC_net_1), .B(controlReg1[3]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[3] ), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] )
        , .Y(), .FCO(\baud_cntr_cry[3] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI3TDS5[2]  (.A(
        VCC_net_1), .B(controlReg1[2]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[2] ), .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] )
        , .Y(), .FCO(\baud_cntr_cry[2] ));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[0] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIB25KC[6]  (.A(
        VCC_net_1), .B(controlReg1[6]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[6] ), .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] )
        , .Y(), .FCO(\baud_cntr_cry[6] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIJB989[4]  (.A(
        VCC_net_1), .B(controlReg1[4]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[4] ), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] )
        , .Y(), .FCO(\baud_cntr_cry[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIU8G64[1]  (.A(
        VCC_net_1), .B(controlReg1[1]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[1] ), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] )
        , .Y(), .FCO(\baud_cntr_cry[1] ));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIMV4OH[9]  (.A(
        VCC_net_1), .B(controlReg2[4]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[9] ), .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] )
        , .Y(), .FCO(\baud_cntr_cry[9] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[6] ));
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        xmit_clock));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNIQ6LQ  (.A(baud_cntr8_8)
        , .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(baud_cntr8_7), .FCI(
        VCC_net_1), .S(), .Y(baud_cntr8_1_RNIQ6LQ_Y), .FCO(
        baud_cntr_cry_cy));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIU57UA[5]  (.A(
        VCC_net_1), .B(controlReg1[5]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[5] ), .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] )
        , .Y(), .FCO(\baud_cntr_cry[5] ));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h44700) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(controlReg2[7]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[12] ), .FCI(\baud_cntr_cry[11] ), .S(
        \baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[1]_net_1 ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI7V31G[8]  (.A(
        VCC_net_1), .B(controlReg2[3]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[8] ), .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] )
        , .Y(), .FCO(\baud_cntr_cry[8] ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[2] ));
    CFG2 #( .INIT(4'h8) )  xmit_pulse_inst_1 (.A(baud_clock), .B(
        xmit_clock), .Y(xmit_pulse));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIEJC2J[10]  (.A(
        VCC_net_1), .B(controlReg2[5]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[10] ), .FCI(\baud_cntr_cry[9] ), .S(
        \baud_cntr_s[10] ), .Y(), .FCO(\baud_cntr_cry[10] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    
endmodule


module mss_sb_CoreUARTapb_2_0_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte_in,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_rx_1
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte_in;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_rx_1;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte_in[7], rx_byte_in[6], 
        rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], 
        rx_byte_in[1], rx_byte_in[0]}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_rx_1), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_ctrl_128_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_2369_i_0,
       N_2370_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_2369_i_0;
input  N_2370_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_empty_rx;
output fifo_full_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[1]_net_1 , VCC_net_1, 
        un1_counter_cry_1_0_S_0, GND_net_1, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_0, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S_0, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_0, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_0, \counter[6]_net_1 , 
        un1_counter_s_6_S_0, \counter[0]_net_1 , un1_counter_cry_0_Y, 
        \data_out_0[0] , \data_out_0[1] , \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \wr_pointer[1]_net_1 , 
        \wr_pointer_s[1] , \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_131_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_132_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_4_net_1, empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_132_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIG41E (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_2_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[2]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_1), 
        .S(un1_counter_cry_2_0_S_0), .Y(), .FCO(un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(N_2369_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_4_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[4]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_3), 
        .S(un1_counter_cry_4_0_S_0), .Y(), .FCO(un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_131_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_131 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_131_FCO));
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_3_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[3]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_2), 
        .S(un1_counter_cry_3_0_S_0), .Y(), .FCO(un1_counter_cry_3));
    ARI1 #( .INIT(20'h56699) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(GND_net_1), .S(), .Y(
        un1_counter_cry_0_Y), .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[2]_net_1 ), .D(\counter[1]_net_1 ), 
        .Y(fifo_empty_rx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_2370_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_1_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_0), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_132 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_132_FCO));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[1]));
    CFG4 #( .INIT(16'h8000) )  full (.A(\counter[0]_net_1 ), .B(
        full_4_net_1), .C(\counter[2]_net_1 ), .D(\counter[1]_net_1 ), 
        .Y(fifo_full_rx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_5_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[5]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_4), 
        .S(un1_counter_cry_5_0_S_0), .Y(), .FCO(un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_0_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte_in({
        rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], 
        rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_rx_1(fifo_write_rx_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(
        \counter[6]_net_1 ), .FCI(un1_counter_cry_5), .S(
        un1_counter_s_6_S_0), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_256x8_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_2369_i_0,
       N_2370_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_2369_i_0;
input  N_2370_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_empty_rx;
output fifo_full_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_0_fifo_ctrl_128_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_byte_in({rx_byte_in[7], 
        rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], 
        rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_2369_i_0(N_2369_i_0), .N_2370_i_0(
        N_2370_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1), .fifo_empty_rx(
        fifo_empty_rx), .fifo_full_rx(fifo_full_rx));
    
endmodule


module mss_sb_CoreUARTapb_2_0_COREUART_1s_1s_0s_15s_0s(
       CoreAPB3_0_APBmslave0_PWDATA,
       data_out,
       controlReg1,
       controlReg2,
       rx_dout_reg_5,
       rx_dout_reg_6,
       rx_dout_reg_7,
       rx_byte_7,
       rx_byte_6,
       rx_byte_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreUARTapb_2_0_OVERFLOW,
       CoreUARTapb_2_0_RXRDY,
       un1_WEn_1,
       CoreAPB3_0_APBmslave2_PSELx,
       un1_WEn_0,
       CoreUARTapb_2_0_PARITY_ERR,
       un1_OEn_2,
       un1_OEn_1,
       BT_RX_c,
       CoreUARTapb_2_0_TXRDY,
       BT_TX_c,
       CoreUARTapb_2_0_FRAMING_ERR
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [4:0] data_out;
input  [7:0] controlReg1;
input  [7:0] controlReg2;
output rx_dout_reg_5;
output rx_dout_reg_6;
output rx_dout_reg_7;
output rx_byte_7;
output rx_byte_6;
output rx_byte_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output CoreUARTapb_2_0_OVERFLOW;
output CoreUARTapb_2_0_RXRDY;
input  un1_WEn_1;
input  CoreAPB3_0_APBmslave2_PSELx;
input  un1_WEn_0;
output CoreUARTapb_2_0_PARITY_ERR;
input  un1_OEn_2;
input  un1_OEn_1;
output BT_RX_c;
output CoreUARTapb_2_0_TXRDY;
input  BT_TX_c;
output CoreUARTapb_2_0_FRAMING_ERR;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, 
        \rx_dout_reg[3]_net_1 , VCC_net_1, \rx_dout[3] , 
        rx_dout_reg4_i_0, GND_net_1, \rx_dout_reg[4]_net_1 , 
        \rx_dout[4] , \rx_dout[5] , \rx_dout[6] , \rx_dout[7] , 
        \tx_hold_reg[0]_net_1 , tx_hold_reg5, \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[4]_net_1 , \tx_hold_reg[5]_net_1 , 
        \tx_hold_reg[6]_net_1 , \tx_hold_reg[7]_net_1 , 
        \rx_dout_reg[0]_net_1 , \rx_dout[0] , \rx_dout_reg[1]_net_1 , 
        \rx_dout[1] , \rx_dout_reg[2]_net_1 , \rx_dout[2] , 
        \rx_state[0]_net_1 , \rx_state_ns[0] , \rx_state[1]_net_1 , 
        N_143_i, rx_dout_reg4, rx_dout_reg_empty_1_sqmuxa_i_0, 
        overflow_reg5_net_1, un1_clear_overflow_net_1, RXRDY5, 
        clear_parity_reg_net_1, clear_parity_reg0, clear_parity_en, 
        fifo_write_tx_net_1, tx_hold_reg5_i_0, fifo_empty_rx, 
        N_2369_i_0, fifo_full_rx, fifo_write, N_2370_i_0, \rx_byte[3] , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[7]_net_1 , 
        \rx_byte_in[6]_net_1 , \rx_byte_in[5]_net_1 , \rx_byte[4] , 
        \rx_byte_in[4]_net_1 , \rx_byte[2] , \rx_byte_in[2]_net_1 , 
        \rx_byte[1] , \rx_byte_in[1]_net_1 , \rx_byte[0] , 
        \rx_byte_in[0]_net_1 , stop_strobe, \rx_state_0[1] , 
        \rx_state_0[0] , fifo_write_rx_1_net_1, fifo_read_rx_0_sqmuxa, 
        xmit_clock, baud_clock, xmit_pulse, \tx_dout_reg[0] , 
        \tx_dout_reg[1] , \tx_dout_reg[2] , \tx_dout_reg[3] , 
        \tx_dout_reg[4] , \tx_dout_reg[5] , \tx_dout_reg[6] , 
        \tx_dout_reg[7] , fifo_read_tx, fifo_read_tx_i_0, 
        fifo_full_tx_i_0, fifo_empty_tx;
    
    SLE \tx_hold_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  overflow_reg5 (.A(fifo_full_rx), .B(
        fifo_write), .Y(overflow_reg5_net_1));
    CFG3 #( .INIT(8'h01) )  fifo_write_rx_1_i (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(N_2370_i_0));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[0]_net_1 ));
    CFG4 #( .INIT(16'hFFFB) )  fifo_read_rx_0_sqmuxa_0_a2_i (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(N_2369_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_143_i));
    CFG3 #( .INIT(8'hFE) )  fifo_write_rx_1 (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(fifo_write_rx_1_net_1));
    mss_sb_CoreUARTapb_2_0_Rx_async_1s_0s_1s_2s make_RX (.rx_byte({
        rx_byte_7, rx_byte_6, rx_byte_5, \rx_byte[4] , \rx_byte[3] , 
        \rx_byte[2] , \rx_byte[1] , \rx_byte[0] }), .rx_state({
        \rx_state_0[1] , \rx_state_0[0] }), .controlReg2({
        controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .clear_parity_reg(clear_parity_reg_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .BT_TX_c(BT_TX_c)
        , .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR), 
        .stop_strobe(stop_strobe), .CoreUARTapb_2_0_FRAMING_ERR(
        CoreUARTapb_2_0_FRAMING_ERR), .clear_parity_en(clear_parity_en)
        , .fifo_write(fifo_write));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[1]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[1] ), .Y(
        \rx_byte_in[1]_net_1 ));
    SLE \tx_hold_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[3]_net_1 ));
    mss_sb_CoreUARTapb_2_0_fifo_256x8 \genblk2.tx_fifo  (.tx_dout_reg({
        \tx_dout_reg[7] , \tx_dout_reg[6] , \tx_dout_reg[5] , 
        \tx_dout_reg[4] , \tx_dout_reg[3] , \tx_dout_reg[2] , 
        \tx_dout_reg[1] , \tx_dout_reg[0] }), .tx_hold_reg({
        \tx_hold_reg[7]_net_1 , \tx_hold_reg[6]_net_1 , 
        \tx_hold_reg[5]_net_1 , \tx_hold_reg[4]_net_1 , 
        \tx_hold_reg[3]_net_1 , \tx_hold_reg[2]_net_1 , 
        \tx_hold_reg[1]_net_1 , \tx_hold_reg[0]_net_1 }), 
        .fifo_write_tx(fifo_write_tx_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[3]  (.A(\rx_byte[3] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[3]_net_1 ), .Y(
        data_out[3]));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE clear_framing_error_reg0 (.D(clear_parity_en), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(clear_parity_reg0));
    SLE \tx_hold_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(GL0_INST), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[5]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_5), .Y(
        \rx_byte_in[5]_net_1 ));
    CFG4 #( .INIT(16'hEEEF) )  \genblk1.RXRDY5  (.A(
        rx_dout_reg_empty_net_1), .B(stop_strobe), .C(\rx_state_0[1] ), 
        .D(\rx_state_0[0] ), .Y(RXRDY5));
    CFG4 #( .INIT(16'h0004) )  fifo_read_rx_0_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(
        fifo_read_rx_0_sqmuxa));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[4]  (.A(\rx_byte[4] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[4]_net_1 ), .Y(
        data_out[4]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[2]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[2] ), .Y(
        \rx_byte_in[2]_net_1 ));
    mss_sb_CoreUARTapb_2_0_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s make_TX (
        .tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .controlReg2({controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .xmit_pulse(
        xmit_pulse), .BT_RX_c(BT_RX_c), .CoreUARTapb_2_0_TXRDY(
        CoreUARTapb_2_0_TXRDY), .fifo_full_tx_i_0(fifo_full_tx_i_0), 
        .xmit_clock(xmit_clock), .baud_clock(baud_clock), 
        .fifo_empty_tx(fifo_empty_tx));
    SLE \tx_hold_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[6]_net_1 ));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[4]_net_1 ));
    mss_sb_CoreUARTapb_2_0_Clock_gen_0s make_CLOCK_GEN (.controlReg1({
        controlReg1[7], controlReg1[6], controlReg1[5], controlReg1[4], 
        controlReg1[3], controlReg1[2], controlReg1[1], controlReg1[0]})
        , .controlReg2({controlReg2[7], controlReg2[6], controlReg2[5], 
        controlReg2[4], controlReg2[3]}), .xmit_clock(xmit_clock), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .xmit_pulse(
        xmit_pulse));
    SLE \rx_state[1]  (.D(N_143_i), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_7));
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hECCC) )  un1_clear_overflow (.A(un1_OEn_2), .B(
        overflow_reg5_net_1), .C(CoreAPB3_0_APBmslave2_PSELx), .D(
        un1_OEn_1), .Y(un1_clear_overflow_net_1));
    SLE clear_parity_reg (.D(clear_parity_reg0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_reg_net_1));
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_5));
    SLE overflow_reg (.D(overflow_reg5_net_1), .CLK(GL0_INST), .EN(
        un1_clear_overflow_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_0_OVERFLOW));
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[0]  (.A(\rx_byte[0] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[0]_net_1 ), .Y(
        data_out[0]));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[2]  (.A(\rx_byte[2] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[2]_net_1 ), .Y(
        data_out[2]));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_6));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \tx_hold_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[7]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(GL0_INST), 
        .EN(RXRDY5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_0_RXRDY));
    mss_sb_CoreUARTapb_2_0_fifo_256x8_0 \genblk3.rx_fifo  (.rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_byte_in({\rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte_in[4]_net_1 , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[1]_net_1 , \rx_byte_in[0]_net_1 }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_2369_i_0(N_2369_i_0), .N_2370_i_0(
        N_2370_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1_net_1), .fifo_empty_rx(
        fifo_empty_rx), .fifo_full_rx(fifo_full_rx));
    SLE \tx_hold_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[3]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \reg_write.tx_hold_reg5_i_0  (.A(un1_WEn_1)
        , .B(CoreAPB3_0_APBmslave2_PSELx), .C(un1_WEn_0), .Y(
        tx_hold_reg5_i_0));
    SLE fifo_write_tx (.D(tx_hold_reg5_i_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_write_tx_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[6]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_6), .Y(
        \rx_byte_in[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[1]  (.A(\rx_byte[1] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[1]_net_1 ), .Y(
        data_out[1]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[7]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_7), .Y(
        \rx_byte_in[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[3]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[3] ), .Y(
        \rx_byte_in[3]_net_1 ));
    SLE \tx_hold_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hB333) )  rx_dout_reg_empty_1_sqmuxa_i (.A(
        un1_OEn_2), .B(rx_dout_reg4), .C(CoreAPB3_0_APBmslave2_PSELx), 
        .D(un1_OEn_1), .Y(rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[4]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[4] ), .Y(
        \rx_byte_in[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[0]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[0] ), .Y(
        \rx_byte_in[0]_net_1 ));
    SLE \tx_hold_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \reg_write.tx_hold_reg5  (.A(un1_WEn_1), 
        .B(CoreAPB3_0_APBmslave2_PSELx), .C(un1_WEn_0), .Y(
        tx_hold_reg5));
    
endmodule


module 
        mss_sb_CoreUARTapb_2_0_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s(
        
       CoreAPB3_0_APBmslave0_PWDATA,
       CoreAPB3_0_APBmslave2_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       un1_OEn_2,
       controlReg24_3,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       un1_OEn_1,
       controlReg24_0,
       controlReg14_3,
       controlReg14_0,
       CoreUARTapb_2_0_PARITY_ERR,
       N_97_1,
       CoreAPB3_0_APBmslave2_PSELx,
       psh_negedge_reg_1_sqmuxa_3_2,
       CoreUARTapb_2_0_FRAMING_ERR,
       CoreUARTapb_2_0_OVERFLOW,
       CoreUARTapb_2_0_RXRDY,
       CoreUARTapb_2_0_TXRDY,
       un1_WEn_1,
       un1_WEn_0,
       BT_RX_c,
       BT_TX_c
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [7:0] CoreAPB3_0_APBmslave2_PRDATA;
input  [4:2] CoreAPB3_0_APBmslave0_PADDR;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output un1_OEn_2;
output controlReg24_3;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
output un1_OEn_1;
output controlReg24_0;
input  controlReg14_3;
output controlReg14_0;
output CoreUARTapb_2_0_PARITY_ERR;
input  N_97_1;
input  CoreAPB3_0_APBmslave2_PSELx;
input  psh_negedge_reg_1_sqmuxa_3_2;
output CoreUARTapb_2_0_FRAMING_ERR;
output CoreUARTapb_2_0_OVERFLOW;
output CoreUARTapb_2_0_RXRDY;
output CoreUARTapb_2_0_TXRDY;
input  un1_WEn_1;
input  un1_WEn_0;
output BT_RX_c;
input  BT_TX_c;

    wire \controlReg1[4]_net_1 , VCC_net_1, controlReg14, GND_net_1, 
        \controlReg1[5]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[7]_net_1 , \NxtPrdata[5] , un1_NxtPrdata23_i_0, 
        \NxtPrdata[6] , \NxtPrdata[7] , \controlReg2[0]_net_1 , 
        controlReg24, \controlReg2[1]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[7]_net_1 , \controlReg1[0]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[3]_net_1 , \NxtPrdata[0] , \NxtPrdata[1] , 
        \NxtPrdata[2] , \NxtPrdata[3] , \NxtPrdata[4] , 
        \NxtPrdata_5_bm[0]_net_1 , \NxtPrdata_5_am[0]_net_1 , 
        \NxtPrdata_5_bm[1]_net_1 , \NxtPrdata_5_am[1]_net_1 , 
        \NxtPrdata_5_bm_0[3] , \NxtPrdata_5_am_0[3] , 
        \NxtPrdata_5_bm_0[4] , \NxtPrdata_5_am_0[4] , 
        \NxtPrdata_5_bm[2]_net_1 , \NxtPrdata_5_am[2]_net_1 , 
        \NxtPrdata_5_bm_0[5] , \NxtPrdata_5_am_0[5] , 
        \NxtPrdata_5_bm_0[7] , \NxtPrdata_5_am_0[7] , 
        \NxtPrdata_5_bm_0[6] , \NxtPrdata_5_am_0[6] , \rx_dout_reg[6] , 
        \rx_byte[6] , \rx_dout_reg[7] , \rx_byte[7] , \rx_dout_reg[5] , 
        \rx_byte[5] , \data_out[2] , \data_out[4] , \data_out[3] , 
        \data_out[1] , \data_out[0] ;
    
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[4]  (.A(
        CoreUARTapb_2_0_FRAMING_ERR), .B(\data_out[4] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[4] ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .C(controlReg24_3), .Y(
        controlReg24_0));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[5]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[5] ), 
        .D(\rx_byte[5] ), .Y(\NxtPrdata_5_am_0[5] ));
    SLE \controlReg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[5]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[0]  (.A(
        CoreUARTapb_2_0_TXRDY), .B(\data_out[0] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[0]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[2]  (.A(
        \controlReg2[2]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[2]_net_1 ), .Y(\NxtPrdata_5_bm[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \p_CtrlReg2Seq.controlReg24_3  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(controlReg24_3));
    SLE \controlReg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[7]_net_1 ));
    SLE \iPRDATA[1]  (.D(\NxtPrdata[1] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[1]));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[6]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[6] ), 
        .D(\rx_byte[6] ), .Y(\NxtPrdata_5_am_0[6] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[7]  (.A(
        \controlReg2[7]_net_1 ), .B(\controlReg1[7]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[7] ));
    SLE \controlReg2[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[4]_net_1 ));
    SLE \iPRDATA[4]  (.D(\NxtPrdata[4] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[4]));
    VCC VCC (.Y(VCC_net_1));
    SLE \iPRDATA[3]  (.D(\NxtPrdata[3] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[3]));
    SLE \controlReg2[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[6]_net_1 ));
    SLE \controlReg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg1Seq.controlReg14  (.A(
        CoreAPB3_0_APBmslave2_PSELx), .B(CoreAPB3_0_APBmslave0_PENABLE)
        , .C(controlReg14_0), .Y(controlReg14));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[4]  (.A(
        \controlReg2[4]_net_1 ), .B(\controlReg1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[4] ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg1Seq.controlReg14_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .C(controlReg14_3), .Y(
        controlReg14_0));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[3]  (.A(
        CoreUARTapb_2_0_OVERFLOW), .B(\data_out[3] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[3] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[5]  (.A(
        \controlReg2[5]_net_1 ), .B(\controlReg1[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[5] ));
    CFG2 #( .INIT(4'h4) )  un1_OEn_2_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(un1_OEn_2));
    CFG3 #( .INIT(8'h02) )  un1_OEn_1_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PENABLE), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PWRITE), .Y(un1_OEn_1));
    SLE \controlReg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[0]  (.A(
        \controlReg2[0]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[0]_net_1 ), .Y(\NxtPrdata_5_bm[0]_net_1 ));
    SLE \controlReg2[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[3]_net_1 ));
    SLE \controlReg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[2]_net_1 ));
    SLE \controlReg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[4]_net_1 ));
    SLE \iPRDATA[5]  (.D(\NxtPrdata[5] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[5]));
    SLE \iPRDATA[7]  (.D(\NxtPrdata[7] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[7]));
    SLE \controlReg2[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[1]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[6]  (.A(
        \controlReg2[6]_net_1 ), .B(\controlReg1[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[6] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[4] ), .C(
        \NxtPrdata_5_am_0[4] ), .Y(\NxtPrdata[4] ));
    SLE \controlReg2[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[7]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24  (.A(
        CoreAPB3_0_APBmslave2_PSELx), .B(CoreAPB3_0_APBmslave0_PENABLE)
        , .C(controlReg24_0), .Y(controlReg24));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[1]_net_1 ), 
        .C(\NxtPrdata_5_am[1]_net_1 ), .Y(\NxtPrdata[1] ));
    SLE \iPRDATA[2]  (.D(\NxtPrdata[2] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[2]));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[0]_net_1 ), 
        .C(\NxtPrdata_5_am[0]_net_1 ), .Y(\NxtPrdata[0] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[3] ), .C(
        \NxtPrdata_5_am_0[3] ), .Y(\NxtPrdata[3] ));
    SLE \controlReg2[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[5]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[3]  (.A(
        \controlReg2[3]_net_1 ), .B(\controlReg1[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[3] ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[1]  (.A(
        CoreUARTapb_2_0_RXRDY), .B(\data_out[1] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[1]_net_1 ));
    SLE \controlReg2[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[2]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  un1_NxtPrdata23_i (.A(
        CoreAPB3_0_APBmslave0_PWRITE), .B(
        CoreAPB3_0_APBmslave0_PENABLE), .C(
        psh_negedge_reg_1_sqmuxa_3_2), .D(CoreAPB3_0_APBmslave2_PSELx), 
        .Y(un1_NxtPrdata23_i_0));
    SLE \iPRDATA[6]  (.D(\NxtPrdata[6] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[6]));
    SLE \iPRDATA[0]  (.D(\NxtPrdata[0] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave2_PRDATA[0]));
    mss_sb_CoreUARTapb_2_0_COREUART_1s_1s_0s_15s_0s uUART (
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .data_out({\data_out[4] , 
        \data_out[3] , \data_out[2] , \data_out[1] , \data_out[0] }), 
        .controlReg1({\controlReg1[7]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[5]_net_1 , \controlReg1[4]_net_1 , 
        \controlReg1[3]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[0]_net_1 }), .controlReg2({
        \controlReg2[7]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[1]_net_1 , \controlReg2[0]_net_1 }), 
        .rx_dout_reg_5(\rx_dout_reg[5] ), .rx_dout_reg_6(
        \rx_dout_reg[6] ), .rx_dout_reg_7(\rx_dout_reg[7] ), 
        .rx_byte_7(\rx_byte[7] ), .rx_byte_6(\rx_byte[6] ), .rx_byte_5(
        \rx_byte[5] ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreUARTapb_2_0_OVERFLOW(CoreUARTapb_2_0_OVERFLOW), 
        .CoreUARTapb_2_0_RXRDY(CoreUARTapb_2_0_RXRDY), .un1_WEn_1(
        un1_WEn_1), .CoreAPB3_0_APBmslave2_PSELx(
        CoreAPB3_0_APBmslave2_PSELx), .un1_WEn_0(un1_WEn_0), 
        .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR), 
        .un1_OEn_2(un1_OEn_2), .un1_OEn_1(un1_OEn_1), .BT_RX_c(BT_RX_c)
        , .CoreUARTapb_2_0_TXRDY(CoreUARTapb_2_0_TXRDY), .BT_TX_c(
        BT_TX_c), .CoreUARTapb_2_0_FRAMING_ERR(
        CoreUARTapb_2_0_FRAMING_ERR));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[7] ), .C(
        \NxtPrdata_5_am_0[7] ), .Y(\NxtPrdata[7] ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[2]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\data_out[2] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[2]_net_1 ));
    SLE \controlReg2[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[0]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[2]_net_1 ), 
        .C(\NxtPrdata_5_am[2]_net_1 ), .Y(\NxtPrdata[2] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[6] ), .C(
        \NxtPrdata_5_am_0[6] ), .Y(\NxtPrdata[6] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[7]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[7] ), 
        .D(\rx_byte[7] ), .Y(\NxtPrdata_5_am_0[7] ));
    SLE \controlReg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[1]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[1]  (.A(
        \controlReg2[1]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[1]_net_1 ), .Y(\NxtPrdata_5_bm[1]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[5] ), .C(
        \NxtPrdata_5_am_0[5] ), .Y(\NxtPrdata[5] ));
    SLE \controlReg1[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[0]_net_1 ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Rx_async_1s_0s_1s_2s(
       rx_byte,
       controlReg2,
       clear_parity_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       GPS_TX_c,
       CoreUARTapb_2_1_PARITY_ERR,
       stop_strobe,
       CoreUARTapb_2_1_FRAMING_ERR,
       clear_parity_en,
       fifo_write,
       rx_idle
    );
output [7:0] rx_byte;
input  [2:0] controlReg2;
input  clear_parity_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  baud_clock;
input  GPS_TX_c;
output CoreUARTapb_2_1_PARITY_ERR;
output stop_strobe;
output CoreUARTapb_2_1_FRAMING_ERR;
output clear_parity_en;
output fifo_write;
output rx_idle;

    wire clear_parity_reg_i_0, \rx_bit_cnt[0]_net_1 , VCC_net_1, 
        N_318_i_0, GND_net_1, \rx_bit_cnt[1]_net_1 , N_319_i_0, 
        \rx_bit_cnt[2]_net_1 , N_320_i_0, \rx_bit_cnt[3]_net_1 , 
        N_321_i_0, \samples[1]_net_1 , \samples[2]_net_1 , 
        \rx_shift[0]_net_1 , \rx_shift_11[0] , 
        un1_samples7_1_0_0_net_1, \rx_shift[1]_net_1 , 
        \rx_shift_11[1] , \rx_shift[2]_net_1 , \rx_shift_11[2] , 
        \rx_shift[3]_net_1 , \rx_shift_11[3] , \rx_shift[4]_net_1 , 
        \rx_shift_11[4] , \rx_shift[5]_net_1 , \rx_shift_11[5] , 
        \rx_shift[6]_net_1 , N_69_i_0, \rx_shift[7]_net_1 , 
        \rx_shift_11[7] , \rx_shift[8]_net_1 , N_71_i_0, 
        \receive_count[0]_net_1 , N_322_i_0, \receive_count[1]_net_1 , 
        N_323_i_0, \receive_count[2]_net_1 , N_324_i_0, 
        \receive_count[3]_net_1 , N_325_i_0, clear_parity_en_9, 
        N_67_i_0, \samples[0]_net_1 , N_310, parity_err_1_sqmuxa_i_0, 
        rx_parity_calc_net_1, N_326_i_0, framing_error_int_net_1, 
        framing_error_int_0_sqmuxa, framing_error_int_2_sqmuxa, 
        framing_error_1_sqmuxa_i_0, \rx_state[1]_net_1 , N_233_i_0, 
        \rx_state[0]_net_1 , \rx_state_ns[0] , clear_parity_en_9_i_0, 
        N_111, N_168, N_172, un1_parity_err_0_sqmuxa_2_1_0_net_1, 
        un1_parity_err_0_sqmuxa_2_1_net_1, rx_state19_li, N_130, N_243, 
        N_112, N_242, framing_error_int_0_sqmuxa_0_a2_2_net_1, N_108, 
        rx_state19_NE_1, N_173, N_118, N_272, un1_parity_err31_1_net_1, 
        N_149, N_116;
    
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[2]_net_1 ));
    CFG4 #( .INIT(16'hE800) )  \rcv_cnt.receive_count_3_i_a2[0]  (.A(
        \samples[0]_net_1 ), .B(\samples[1]_net_1 ), .C(
        \samples[2]_net_1 ), .D(rx_idle), .Y(N_172));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[0]));
    CFG4 #( .INIT(16'h0004) )  \rcv_cnt.receive_count_3_i_a2_0[3]  (.A(
        \receive_count[0]_net_1 ), .B(rx_idle), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_272));
    SLE \receive_count[1]  (.D(N_323_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[1]_net_1 ));
    SLE \rx_shift[7]  (.D(\rx_shift_11[7] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[7]_net_1 ));
    CFG4 #( .INIT(16'h0096) )  
        \make_parity_err.parity_err_12_iv_0_111_a2  (.A(controlReg2[2])
        , .B(rx_parity_calc_net_1), .C(N_118), .D(clear_parity_reg), 
        .Y(N_310));
    CFG3 #( .INIT(8'h08) )  framing_error_int_0_sqmuxa_0_a2_2 (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(
        framing_error_int_0_sqmuxa_0_a2_2_net_1));
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[0]_net_1 ));
    CFG3 #( .INIT(8'h40) )  
        \receive_full_indicator.clear_parity_en_9_0_a3  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9));
    CFG3 #( .INIT(8'h10) )  un1_samples7_1_0_0_a2 (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .C(baud_clock), 
        .Y(N_168));
    CFG2 #( .INIT(4'hE) )  \receive_shift.rx_shift_11_i_o2[6]  (.A(
        controlReg2[1]), .B(controlReg2[0]), .Y(N_112));
    CFG1 #( .INIT(2'h1) )  framing_error_RNO (.A(clear_parity_reg), .Y(
        clear_parity_reg_i_0));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[0]  (.A(rx_idle), 
        .B(\rx_shift[1]_net_1 ), .Y(\rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(N_325_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hDF) )  un1_samples7_1_0_0_o2 (.A(baud_clock), .B(
        N_108), .C(\receive_count[3]_net_1 ), .Y(N_111));
    CFG2 #( .INIT(4'h1) )  \rx_state_ns_0_a3_0_3_0_a2[0]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(rx_idle));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[4]));
    CFG4 #( .INIT(16'h333B) )  un1_samples7_1_0_0 (.A(baud_clock), .B(
        N_111), .C(\rx_state[1]_net_1 ), .D(\rx_state[0]_net_1 ), .Y(
        un1_samples7_1_0_0_net_1));
    CFG3 #( .INIT(8'h7F) )  un1_parity_err31_1 (.A(controlReg2[1]), .B(
        baud_clock), .C(un1_parity_err_0_sqmuxa_2_1_net_1), .Y(
        un1_parity_err31_1_net_1));
    SLE rx_parity_calc (.D(N_326_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_parity_calc_net_1));
    SLE \rx_bit_cnt[2]  (.D(N_320_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[2]_net_1 ));
    SLE \rx_bit_cnt[1]  (.D(N_319_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[1]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  \rcv_cnt.receive_count_3_i_a2_0[0]  (.A(
        \receive_count[1]_net_1 ), .B(\receive_count[2]_net_1 ), .C(
        rx_idle), .D(\receive_count[3]_net_1 ), .Y(N_173));
    CFG3 #( .INIT(8'h7F) )  \rcv_cnt.receive_count_3_i_o2[2]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(N_108));
    CFG3 #( .INIT(8'h21) )  rx_parity_calc_RNO (.A(
        rx_parity_calc_net_1), .B(\rx_state[1]_net_1 ), .C(N_149), .Y(
        N_326_i_0));
    CFG3 #( .INIT(8'hDF) )  \receive_shift.rx_bit_cnt_4_i_o2[1]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(N_111), .C(\rx_bit_cnt[1]_net_1 ), 
        .Y(N_116));
    CFG4 #( .INIT(16'h00E4) )  \receive_shift.rx_shift_11[7]  (.A(
        N_243), .B(N_242), .C(N_118), .D(rx_idle), .Y(\rx_shift_11[7] )
        );
    CFG3 #( .INIT(8'h09) )  \rx_bit_cnt_RNO[0]  (.A(N_111), .B(
        \rx_bit_cnt[0]_net_1 ), .C(N_168), .Y(N_318_i_0));
    CFG4 #( .INIT(16'h1230) )  \receive_count_RNO[2]  (.A(
        \receive_count[0]_net_1 ), .B(N_172), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_324_i_0));
    CFG3 #( .INIT(8'hAC) )  \receive_shift.rx_shift_9_0[7]  (.A(
        \rx_shift[8]_net_1 ), .B(\rx_shift[7]_net_1 ), .C(
        controlReg2[1]), .Y(N_242));
    CFG4 #( .INIT(16'hFDBF) )  \rcv_sm.rx_state19_NE_1  (.A(
        \rx_bit_cnt[1]_net_1 ), .B(N_112), .C(\rx_bit_cnt[3]_net_1 ), 
        .D(\rx_bit_cnt[2]_net_1 ), .Y(rx_state19_NE_1));
    SLE stop_strobe_inst_1 (.D(framing_error_int_2_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG4 #( .INIT(16'h0D08) )  \rx_shift_RNO[6]  (.A(N_112), .B(
        \rx_shift[7]_net_1 ), .C(rx_idle), .D(N_118), .Y(N_69_i_0));
    CFG4 #( .INIT(16'h00CE) )  \rx_state_RNO[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .C(
        rx_state19_li), .D(framing_error_int_2_sqmuxa), .Y(N_233_i_0));
    CFG3 #( .INIT(8'h09) )  \rx_bit_cnt_RNO[2]  (.A(N_116), .B(
        \rx_bit_cnt[2]_net_1 ), .C(N_168), .Y(N_320_i_0));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[1]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[2]  (.A(rx_idle), 
        .B(\rx_shift[3]_net_1 ), .Y(\rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(N_324_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[2]_net_1 ));
    SLE clear_parity_en_1 (.D(clear_parity_en_9), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_en));
    CFG4 #( .INIT(16'h4008) )  un1_parity_err_0_sqmuxa_2_1 (.A(
        controlReg2[0]), .B(un1_parity_err_0_sqmuxa_2_1_0_net_1), .C(
        \rx_bit_cnt[1]_net_1 ), .D(\rx_bit_cnt[0]_net_1 ), .Y(
        un1_parity_err_0_sqmuxa_2_1_net_1));
    SLE \rx_state[1]  (.D(N_233_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[6]));
    CFG3 #( .INIT(8'h12) )  \receive_count_RNO[1]  (.A(
        \receive_count[0]_net_1 ), .B(N_172), .C(
        \receive_count[1]_net_1 ), .Y(N_323_i_0));
    GND GND (.Y(GND_net_1));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[3]  (.A(rx_idle), 
        .B(\rx_shift[4]_net_1 ), .Y(\rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(N_67_i_0), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[7]));
    CFG3 #( .INIT(8'hEB) )  \rcv_sm.rx_state19_NE  (.A(rx_state19_NE_1)
        , .B(\rx_bit_cnt[0]_net_1 ), .C(N_243), .Y(rx_state19_li));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[3]));
    CFG4 #( .INIT(16'h0009) )  \receive_count_RNO[3]  (.A(N_108), .B(
        \receive_count[3]_net_1 ), .C(N_172), .D(N_272), .Y(N_325_i_0));
    CFG3 #( .INIT(8'h20) )  \rx_state_ns_i_a3_0_0_a2[1]  (.A(
        \receive_count[3]_net_1 ), .B(N_108), .C(\rx_state[1]_net_1 ), 
        .Y(framing_error_int_2_sqmuxa));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[2]));
    CFG3 #( .INIT(8'h42) )  un1_parity_err_0_sqmuxa_2_1_0 (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(
        \rx_bit_cnt[1]_net_1 ), .Y(un1_parity_err_0_sqmuxa_2_1_0_net_1)
        );
    CFG3 #( .INIT(8'hE8) )  \rx_filtered.m3_0_o2  (.A(
        \samples[1]_net_1 ), .B(\samples[0]_net_1 ), .C(
        \samples[2]_net_1 ), .Y(N_118));
    CFG3 #( .INIT(8'h01) )  \receive_count_RNO[0]  (.A(N_172), .B(
        \receive_count[0]_net_1 ), .C(N_173), .Y(N_322_i_0));
    CFG2 #( .INIT(4'h7) )  \receive_shift.rx_shift_11_i_o2[8]  (.A(
        controlReg2[1]), .B(controlReg2[0]), .Y(N_130));
    SLE parity_err (.D(N_310), .CLK(GL0_INST), .EN(
        parity_err_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_1_PARITY_ERR));
    SLE \rx_shift[6]  (.D(N_69_i_0), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[6]_net_1 ));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[4]  (.A(rx_idle), 
        .B(\rx_shift[5]_net_1 ), .Y(\rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[3]_net_1 ));
    SLE framing_error_int (.D(framing_error_int_0_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(framing_error_int_net_1));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \samples[2]  (.D(GPS_TX_c), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    SLE \receive_count[0]  (.D(N_322_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[5]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[5]  (.A(rx_idle), 
        .B(\rx_shift[6]_net_1 ), .Y(\rx_shift_11[5] ));
    CFG3 #( .INIT(8'hBF) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_i  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9_i_0));
    CFG4 #( .INIT(16'h2000) )  framing_error_int_0_sqmuxa_0_a2 (.A(
        framing_error_int_0_sqmuxa_0_a2_2_net_1), .B(N_118), .C(
        \rx_state[1]_net_1 ), .D(\receive_count[3]_net_1 ), .Y(
        framing_error_int_0_sqmuxa));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[5]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \rx_state_ns_0[0]  (.A(N_272), .B(
        rx_state19_li), .C(\rx_state[0]_net_1 ), .D(
        \receive_count[3]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_bit_cnt[0]  (.D(N_318_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[0]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  framing_error_1_sqmuxa_i (.A(
        framing_error_int_net_1), .B(clear_parity_reg), .C(baud_clock), 
        .Y(framing_error_1_sqmuxa_i_0));
    SLE \rx_shift[8]  (.D(N_71_i_0), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[1]  (.A(rx_idle), 
        .B(\rx_shift[2]_net_1 ), .Y(\rx_shift_11[1] ));
    SLE framing_error (.D(clear_parity_reg_i_0), .CLK(GL0_INST), .EN(
        framing_error_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_1_FRAMING_ERR));
    CFG4 #( .INIT(16'hFF7F) )  \rx_par_calc.rx_parity_calc_4_u_i_o2  (
        .A(controlReg2[1]), .B(\receive_count[3]_net_1 ), .C(N_118), 
        .D(N_108), .Y(N_149));
    CFG4 #( .INIT(16'h3022) )  \rx_shift_RNO[8]  (.A(N_118), .B(
        rx_idle), .C(\rx_shift[8]_net_1 ), .D(N_130), .Y(N_71_i_0));
    CFG2 #( .INIT(4'h6) )  \receive_shift.rx_shift_9_sn_m1  (.A(
        controlReg2[1]), .B(controlReg2[0]), .Y(N_243));
    CFG2 #( .INIT(4'h8) )  \rx_byte_RNO[7]  (.A(controlReg2[0]), .B(
        \rx_shift[7]_net_1 ), .Y(N_67_i_0));
    CFG4 #( .INIT(16'h0A06) )  \rx_bit_cnt_RNO[3]  (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(N_168), 
        .D(N_116), .Y(N_321_i_0));
    CFG4 #( .INIT(16'hCCCE) )  parity_err_1_sqmuxa_i (.A(
        \receive_count[3]_net_1 ), .B(clear_parity_reg), .C(
        un1_parity_err31_1_net_1), .D(N_108), .Y(
        parity_err_1_sqmuxa_i_0));
    SLE \rx_bit_cnt[3]  (.D(N_321_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h0A06) )  \rx_bit_cnt_RNO[1]  (.A(
        \rx_bit_cnt[1]_net_1 ), .B(\rx_bit_cnt[0]_net_1 ), .C(N_168), 
        .D(N_111), .Y(N_319_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_1_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] tx_hold_reg;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), .C_WEN(
        INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), 
        .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_ctrl_128(
       counter,
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_full_tx_i_0
    );
output [6:0] counter;
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_2336_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, VCC_net_1, 
        un1_counter_cry_0_Y_1, GND_net_1, un1_counter_cry_1_0_S_1, 
        un1_counter_cry_2_0_S_1, un1_counter_cry_3_0_S_1, 
        un1_counter_cry_4_0_S_1, un1_counter_cry_5_0_S_1, 
        un1_counter_s_6_S_1, \data_out_0[2] , \data_out_0[3] , 
        \data_out_0[4] , \data_out_0[5] , \data_out_0[6] , 
        \data_out_0[7] , \data_out_0[0] , \data_out_0[1] , 
        \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_125_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_126_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_0_a2_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_126_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[2]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_2_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(counter[2]), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S_1), .Y(), .FCO(
        un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[6]));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_4_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(counter[4]), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S_1), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_125_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[4]));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_126 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_126_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[4]));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[5]));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[5]));
    CFG4 #( .INIT(16'h7FFF) )  full_0_a2_4_RNIKNHS (.A(counter[0]), .B(
        full_0_a2_4_net_1), .C(counter[5]), .D(counter[4]), .Y(
        fifo_full_tx_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_0_a2_4 (.A(counter[6]), .B(
        counter[3]), .C(counter[2]), .D(counter[1]), .Y(
        full_0_a2_4_net_1));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[1]));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[3]));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[6]));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_3_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(counter[3]), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S_1), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(counter[0]), .B(
        fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(un1_counter_cry_0_Y_1), .FCO(
        un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNII4ID (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_2336_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_2336_i_0 (.A(fifo_write_tx), .Y(
        N_2336_i_0_net_1));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_125 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_125_FCO));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_1_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(counter[1]), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_1), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_5_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(counter[5]), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S_1), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_1_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg({
        tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], 
        tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]})
        , .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_tx(fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(counter[6]), .FCI(
        un1_counter_cry_5), .S(un1_counter_s_6_S_1), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        counter[0]));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_256x8(
       counter,
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_full_tx_i_0
    );
output [6:0] counter;
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_1_fifo_ctrl_128 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.counter({counter[6], 
        counter[5], counter[4], counter[3], counter[2], counter[1], 
        counter[0]}), .tx_dout_reg({tx_dout_reg[7], tx_dout_reg[6], 
        tx_dout_reg[5], tx_dout_reg[4], tx_dout_reg[3], tx_dout_reg[2], 
        tx_dout_reg[1], tx_dout_reg[0]}), .tx_hold_reg({tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), 
        .fifo_write_tx(fifo_write_tx), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       counter,
       controlReg2,
       fifo_read_tx,
       fifo_read_tx_i_0,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_110,
       GPS_RX_c,
       CoreUARTapb_2_1_TXRDY,
       fifo_full_tx_i_0,
       xmit_clock,
       baud_clock
    );
input  [7:0] tx_dout_reg;
input  [6:0] counter;
input  [2:0] controlReg2;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_110;
output GPS_RX_c;
output CoreUARTapb_2_1_TXRDY;
input  fifo_full_tx_i_0;
input  xmit_clock;
input  baud_clock;

    wire \tx_byte[4]_net_1 , VCC_net_1, N_123_i_0, GND_net_1, 
        \tx_byte[5]_net_1 , \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_122_i_0, \xmit_bit_sel[2]_net_1 , 
        N_124_i_0, \xmit_bit_sel[3]_net_1 , N_126_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , \tx_byte[2]_net_1 , 
        \tx_byte[3]_net_1 , tx_parity_net_1, N_84_i_0, 
        un1_tx_parity_1_sqmuxa_0_0_net_1, tx_4_iv_i_0, N_81, 
        fifo_read_en0_1_i_a3_i_net_1, \xmit_state[6]_net_1 , N_327_i_0, 
        \xmit_state[0]_net_1 , \xmit_state_ns[0] , 
        \xmit_state[1]_net_1 , \xmit_state[2]_net_1 , 
        \xmit_state_ns[2] , \xmit_state[3]_net_1 , N_112_i_0, 
        \xmit_state[4]_net_1 , \xmit_state_ns[4] , 
        \xmit_state[5]_net_1 , \xmit_state_ns[5] , N_271, 
        tx_2_u_i_m2_am_1_1, tx_2_u_i_m2_am, tx_2_u_i_m2_bm_1_1, 
        tx_2_u_i_m2_bm, N_142, \xmit_state_ns_0_a2_0_4[0]_net_1 , 
        \xmit_state_ns_0_a2_0_5[0]_net_1 , N_114, N_107_i, N_192, 
        N_276, N_165;
    
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(
        tx_2_u_i_m2_bm_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_bm));
    CFG2 #( .INIT(4'h7) )  \xmit_cnt.xmit_bit_sel_3_i_0_o2[2]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        N_114));
    SLE tx_parity (.D(N_84_i_0), .CLK(GL0_INST), .EN(
        un1_tx_parity_1_sqmuxa_0_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_parity_net_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_1_TXRDY));
    CFG4 #( .INIT(16'h8000) )  un1_tx_parity_1_sqmuxa_0_0_a2 (.A(
        \xmit_state[3]_net_1 ), .B(xmit_clock), .C(baud_clock), .D(
        controlReg2[1]), .Y(N_271));
    CFG3 #( .INIT(8'hD8) )  \xmit_sel.tx_2_u_i_m2_ns  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(tx_2_u_i_m2_bm), .C(
        tx_2_u_i_m2_am), .Y(N_142));
    SLE \xmit_state[3]  (.D(N_112_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[3]_net_1 ));
    CFG3 #( .INIT(8'h82) )  \xmit_sel.tx_4_iv_0_a2  (.A(
        \xmit_state[4]_net_1 ), .B(controlReg2[2]), .C(tx_parity_net_1)
        , .Y(N_192));
    CFG4 #( .INIT(16'h0001) )  \xmit_state_ns_0_a2_0_5[0]  (.A(
        counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[0]), 
        .Y(\xmit_state_ns_0_a2_0_5[0]_net_1 ));
    CFG4 #( .INIT(16'h0031) )  \xmit_sel.tx_4_iv_i  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(N_142), 
        .D(N_192), .Y(tx_4_iv_i_0));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[0]_net_1 ));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[4]_net_1 ));
    CFG4 #( .INIT(16'hFFAC) )  \xmit_state_ns_0[5]  (.A(
        \xmit_state[4]_net_1 ), .B(\xmit_state[5]_net_1 ), .C(N_110), 
        .D(N_165), .Y(\xmit_state_ns[5] ));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns_0[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(N_110), 
        .Y(\xmit_state_ns[2] ));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3_0_a2[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[0]_net_1 ), .B(\xmit_bit_sel[1]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_122_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNI2248 (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[5]_net_1 ));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_bm_1_1));
    CFG3 #( .INIT(8'h12) )  tx_parity_RNO (.A(tx_parity_net_1), .B(
        \xmit_state[5]_net_1 ), .C(N_142), .Y(N_84_i_0));
    CFG2 #( .INIT(4'h6) )  \xmit_state_ns_0_x2[4]  (.A(controlReg2[0]), 
        .B(\xmit_bit_sel[0]_net_1 ), .Y(N_107_i));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  \xmit_state_ns_0_a2_0_4[0]  (.A(
        counter[4]), .B(\xmit_state[0]_net_1 ), .C(counter[6]), .D(
        counter[5]), .Y(\xmit_state_ns_0_a2_0_4[0]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \xmit_state_ns_0_a2[5]  (.A(
        \xmit_state[3]_net_1 ), .B(controlReg2[1]), .C(N_276), .D(
        N_110), .Y(N_165));
    CFG3 #( .INIT(8'h4C) )  fifo_read_en0_1_i_a3_i_i (.A(
        \xmit_state_ns_0_a2_0_4[0]_net_1 ), .B(\xmit_state[0]_net_1 ), 
        .C(\xmit_state_ns_0_a2_0_5[0]_net_1 ), .Y(N_327_i_0));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_126_i_0), .CLK(GL0_INST), .EN(N_110), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[3]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns_0[0]  (.A(
        \xmit_state[5]_net_1 ), .B(\xmit_state_ns_0_a2_0_5[0]_net_1 ), 
        .C(\xmit_state_ns_0_a2_0_4[0]_net_1 ), .D(N_110), .Y(
        \xmit_state_ns[0] ));
    SLE \xmit_bit_sel[2]  (.D(N_124_i_0), .CLK(GL0_INST), .EN(N_110), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE tx (.D(tx_4_iv_i_0), .CLK(GL0_INST), .EN(N_81), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(GPS_RX_c));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[3]_net_1 ));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[7]_net_1 ));
    CFG4 #( .INIT(16'hCAEA) )  \xmit_state_RNO[3]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(N_110), 
        .D(N_276), .Y(N_112_i_0));
    CFG3 #( .INIT(8'h84) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_114), 
        .Y(N_124_i_0));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[6]_net_1 ));
    CFG4 #( .INIT(16'h0200) )  \xmit_state_ns_0_a2_1[4]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(N_107_i), .C(
        \xmit_bit_sel[3]_net_1 ), .D(\xmit_bit_sel[2]_net_1 ), .Y(
        N_276));
    CFG2 #( .INIT(4'hE) )  un1_tx_parity_1_sqmuxa_0_0 (.A(N_271), .B(
        \xmit_state[5]_net_1 ), .Y(un1_tx_parity_1_sqmuxa_0_0_net_1));
    SLE \xmit_bit_sel[1]  (.D(N_122_i_0), .CLK(GL0_INST), .EN(N_110), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[1]_net_1 ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[1]_net_1 ));
    CFG4 #( .INIT(16'hAE0C) )  \xmit_state_ns_0[4]  (.A(N_271), .B(
        \xmit_state[4]_net_1 ), .C(N_110), .D(N_276), .Y(
        \xmit_state_ns[4] ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(GL0_INST), 
        .EN(N_110), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[2]_net_1 ));
    SLE fifo_read_en0 (.D(fifo_read_en0_1_i_a3_i_net_1), .CLK(GL0_INST)
        , .EN(N_81), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    CFG2 #( .INIT(4'h8) )  \xmit_state_RNI093E[2]  (.A(N_110), .B(
        \xmit_state[2]_net_1 ), .Y(N_123_i_0));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(GL0_INST), .EN(
        N_123_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[1]_net_1 ));
    SLE \xmit_state[4]  (.D(\xmit_state_ns[4] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[4]_net_1 ));
    CFG4 #( .INIT(16'hC600) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_bit_sel[3]_net_1 ), .C(
        N_114), .D(\xmit_state[3]_net_1 ), .Y(N_126_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_am_1_1));
    SLE \xmit_state[6]  (.D(N_327_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[6]_net_1 ));
    CFG3 #( .INIT(8'hB3) )  fifo_read_en0_1_i_a3_i (.A(
        \xmit_state_ns_0_a2_0_4[0]_net_1 ), .B(\xmit_state[0]_net_1 ), 
        .C(\xmit_state_ns_0_a2_0_5[0]_net_1 ), .Y(
        fifo_read_en0_1_i_a3_i_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_sm.fifo_read_en020_i_a3_i  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(N_110), 
        .D(\xmit_state[6]_net_1 ), .Y(N_81));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(
        tx_2_u_i_m2_am_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_am));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Clock_gen_0s(
       controlReg1,
       controlReg2,
       xmit_clock,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       N_110
    );
input  [7:0] controlReg1;
input  [7:3] controlReg2;
output xmit_clock;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output baud_clock;
output N_110;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNIURC7_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIM2N85[9]  (.A(
        VCC_net_1), .B(controlReg2[4]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[9] ), .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] )
        , .Y(), .FCO(\baud_cntr_cry[9] ));
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[1] ));
    CFG2 #( .INIT(4'h8) )  xmit_pulse_0_o2 (.A(baud_clock), .B(
        xmit_clock), .Y(N_110));
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[3] ));
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[3]_net_1 ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI61172[3]  (.A(
        VCC_net_1), .B(controlReg1[3]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[3] ), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] )
        , .Y(), .FCO(\baud_cntr_cry[3] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIE7M64[7]  (.A(
        VCC_net_1), .B(controlReg1[7]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[7] ), .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] )
        , .Y(), .FCO(\baud_cntr_cry[7] ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[9] ));
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNIURC7_Y), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(baud_clock));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIK58R5[10]  (.A(
        VCC_net_1), .B(controlReg2[5]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[10] ), .FCI(\baud_cntr_cry[9] ), .S(
        \baud_cntr_s[10] ), .Y(), .FCO(\baud_cntr_cry[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI6GR63[5]  (.A(
        VCC_net_1), .B(controlReg1[5]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[5] ), .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] )
        , .Y(), .FCO(\baud_cntr_cry[5] ));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[7] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI1KMN4[8]  (.A(
        VCC_net_1), .B(controlReg2[3]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[8] ), .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] )
        , .Y(), .FCO(\baud_cntr_cry[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIEQ671[1]  (.A(
        VCC_net_1), .B(controlReg1[1]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[1] ), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] )
        , .Y(), .FCO(\baud_cntr_cry[1] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[5] ));
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIKAPD6[11]  (.A(
        VCC_net_1), .B(controlReg2[6]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[11] ), .FCI(\baud_cntr_cry[10] ), .S(
        \baud_cntr_s[11] ), .Y(), .FCO(\baud_cntr_cry[11] ));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNIURC7  (.A(baud_cntr8_8)
        , .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(baud_cntr8_7), .FCI(
        VCC_net_1), .S(), .Y(baud_cntr8_1_RNIURC7_Y), .FCO(
        baud_cntr_cry_cy));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[0] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIPS3N1[2]  (.A(
        VCC_net_1), .B(controlReg1[2]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[2] ), .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] )
        , .Y(), .FCO(\baud_cntr_cry[2] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[6] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI5Q9N[0]  (.A(
        VCC_net_1), .B(controlReg1[0]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[0] ), .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), 
        .Y(), .FCO(\baud_cntr_cry[0] ));
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        xmit_clock));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h44700) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(controlReg2[7]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[12] ), .FCI(\baud_cntr_cry[11] ), .S(
        \baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[1]_net_1 ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIL7UM2[4]  (.A(
        VCC_net_1), .B(controlReg1[4]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[4] ), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] )
        , .Y(), .FCO(\baud_cntr_cry[4] ));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIPQOM3[6]  (.A(
        VCC_net_1), .B(controlReg1[6]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[6] ), .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] )
        , .Y(), .FCO(\baud_cntr_cry[6] ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte_in,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_rx_1
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte_in;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_rx_1;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte_in[7], rx_byte_in[6], 
        rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], 
        rx_byte_in[1], rx_byte_in[0]}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_rx_1), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_ctrl_128_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_2318_i_0,
       N_2319_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_full_rx,
       fifo_empty_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_2318_i_0;
input  N_2319_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_full_rx;
output fifo_empty_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[1]_net_1 , VCC_net_1, 
        un1_counter_cry_1_0_S_2, GND_net_1, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_2, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S_2, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_2, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_2, \counter[6]_net_1 , 
        un1_counter_s_6_S_2, \counter[0]_net_1 , un1_counter_cry_0_Y_2, 
        \data_out_0[0] , \data_out_0[1] , \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \wr_pointer[1]_net_1 , 
        \wr_pointer_s[1] , \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_127_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_128_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_4_net_1, empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_128_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIHD74 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_2_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[2]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_1), 
        .S(un1_counter_cry_2_0_S_2), .Y(), .FCO(un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(N_2318_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_4_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[4]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_3), 
        .S(un1_counter_cry_4_0_S_2), .Y(), .FCO(un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_127_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_3_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[3]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_2), 
        .S(un1_counter_cry_3_0_S_2), .Y(), .FCO(un1_counter_cry_3));
    ARI1 #( .INIT(20'h56699) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(GND_net_1), .S(), .Y(
        un1_counter_cry_0_Y_2), .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[2]_net_1 ), .D(\counter[1]_net_1 ), 
        .Y(fifo_empty_rx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_2319_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_1_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_2), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[1]));
    CFG4 #( .INIT(16'h8000) )  full (.A(\counter[0]_net_1 ), .B(
        full_4_net_1), .C(\counter[2]_net_1 ), .D(\counter[1]_net_1 ), 
        .Y(fifo_full_rx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_5_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[5]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_4), 
        .S(un1_counter_cry_5_0_S_2), .Y(), .FCO(un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_1_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte_in({
        rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], 
        rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_rx_1(fifo_write_rx_1));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_127 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_127_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(
        \counter[6]_net_1 ), .FCI(un1_counter_cry_5), .S(
        un1_counter_s_6_S_2), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_128 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_128_FCO));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_256x8_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_2318_i_0,
       N_2319_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_full_rx,
       fifo_empty_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_2318_i_0;
input  N_2319_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_full_rx;
output fifo_empty_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_1_fifo_ctrl_128_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_byte_in({rx_byte_in[7], 
        rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], 
        rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_2318_i_0(N_2318_i_0), .N_2319_i_0(
        N_2319_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1), .fifo_full_rx(fifo_full_rx), 
        .fifo_empty_rx(fifo_empty_rx));
    
endmodule


module mss_sb_CoreUARTapb_2_1_COREUART_1s_1s_0s_15s_0s(
       CoreAPB3_0_APBmslave0_PWDATA,
       data_out,
       controlReg1,
       controlReg2,
       rx_dout_reg_5,
       rx_dout_reg_6,
       rx_dout_reg_7,
       rx_dout_reg_0,
       rx_dout_reg_1,
       rx_dout_reg_2,
       rx_byte_5,
       rx_byte_0,
       rx_byte_2,
       rx_byte_1,
       rx_byte_6,
       rx_byte_7,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreUARTapb_2_1_OVERFLOW,
       CoreUARTapb_2_1_RXRDY,
       un1_WEn_1,
       CoreAPB3_0_APBmslave3_PSELx,
       un1_WEn_0,
       CoreUARTapb_2_1_PARITY_ERR,
       un1_OEn_2,
       un1_OEn_1,
       GPS_RX_c,
       CoreUARTapb_2_1_TXRDY,
       GPS_TX_c,
       CoreUARTapb_2_1_FRAMING_ERR
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [4:3] data_out;
input  [7:0] controlReg1;
input  [7:0] controlReg2;
output rx_dout_reg_5;
output rx_dout_reg_6;
output rx_dout_reg_7;
output rx_dout_reg_0;
output rx_dout_reg_1;
output rx_dout_reg_2;
output rx_byte_5;
output rx_byte_0;
output rx_byte_2;
output rx_byte_1;
output rx_byte_6;
output rx_byte_7;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output CoreUARTapb_2_1_OVERFLOW;
output CoreUARTapb_2_1_RXRDY;
input  un1_WEn_1;
input  CoreAPB3_0_APBmslave3_PSELx;
input  un1_WEn_0;
output CoreUARTapb_2_1_PARITY_ERR;
input  un1_OEn_2;
input  un1_OEn_1;
output GPS_RX_c;
output CoreUARTapb_2_1_TXRDY;
input  GPS_TX_c;
output CoreUARTapb_2_1_FRAMING_ERR;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, 
        \rx_dout_reg[3]_net_1 , VCC_net_1, \rx_dout[3] , 
        rx_dout_reg4_i_0, GND_net_1, \rx_dout_reg[4]_net_1 , 
        \rx_dout[4] , \rx_dout[5] , \rx_dout[6] , \rx_dout[7] , 
        \tx_hold_reg[0]_net_1 , tx_hold_reg5, \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[4]_net_1 , \tx_hold_reg[5]_net_1 , 
        \tx_hold_reg[6]_net_1 , \tx_hold_reg[7]_net_1 , \rx_dout[0] , 
        \rx_dout[1] , \rx_dout[2] , \rx_state[0]_net_1 , 
        \rx_state_ns[0] , \rx_state[1]_net_1 , N_143_i, rx_dout_reg4, 
        rx_dout_reg_empty_1_sqmuxa_i_0, overflow_reg5_net_1, 
        un1_clear_overflow_0, RXRDY5, clear_parity_reg_net_1, 
        clear_parity_reg0, clear_parity_en, fifo_write_tx_net_1, 
        tx_hold_reg5_i_0, fifo_empty_rx, N_2318_i_0, fifo_full_rx, 
        fifo_write, N_2319_i_0, \rx_byte_in[5]_net_1 , 
        \rx_byte_in[0]_net_1 , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[1]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[7]_net_1 , \rx_byte[4] , \rx_byte_in[4]_net_1 , 
        \rx_byte[3] , \rx_byte_in[3]_net_1 , rx_idle, stop_strobe, 
        fifo_write_rx_1_net_1, fifo_read_rx_0_sqmuxa, xmit_clock, 
        baud_clock, N_110, \tx_dout_reg[0] , \tx_dout_reg[1] , 
        \tx_dout_reg[2] , \tx_dout_reg[3] , \tx_dout_reg[4] , 
        \tx_dout_reg[5] , \tx_dout_reg[6] , \tx_dout_reg[7] , 
        \counter[0] , \counter[1] , \counter[2] , \counter[3] , 
        \counter[4] , \counter[5] , \counter[6] , fifo_read_tx, 
        fifo_read_tx_i_0, fifo_full_tx_i_0;
    
    SLE \tx_hold_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  overflow_reg5 (.A(fifo_full_rx), .B(
        fifo_write), .Y(overflow_reg5_net_1));
    CFG3 #( .INIT(8'h01) )  fifo_write_rx_1_i (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(N_2319_i_0));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_0));
    CFG4 #( .INIT(16'hFFFB) )  fifo_read_rx_0_sqmuxa_0_a2_i (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(N_2318_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_143_i));
    CFG3 #( .INIT(8'hFE) )  fifo_write_rx_1 (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(fifo_write_rx_1_net_1));
    mss_sb_CoreUARTapb_2_1_Rx_async_1s_0s_1s_2s make_RX (.rx_byte({
        rx_byte_7, rx_byte_6, rx_byte_5, \rx_byte[4] , \rx_byte[3] , 
        rx_byte_2, rx_byte_1, rx_byte_0}), .controlReg2({
        controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .clear_parity_reg(clear_parity_reg_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .GPS_TX_c(
        GPS_TX_c), .CoreUARTapb_2_1_PARITY_ERR(
        CoreUARTapb_2_1_PARITY_ERR), .stop_strobe(stop_strobe), 
        .CoreUARTapb_2_1_FRAMING_ERR(CoreUARTapb_2_1_FRAMING_ERR), 
        .clear_parity_en(clear_parity_en), .fifo_write(fifo_write), 
        .rx_idle(rx_idle));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[1]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_1), .Y(
        \rx_byte_in[1]_net_1 ));
    SLE \tx_hold_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[3]_net_1 ));
    mss_sb_CoreUARTapb_2_1_fifo_256x8 \genblk2.tx_fifo  (.counter({
        \counter[6] , \counter[5] , \counter[4] , \counter[3] , 
        \counter[2] , \counter[1] , \counter[0] }), .tx_dout_reg({
        \tx_dout_reg[7] , \tx_dout_reg[6] , \tx_dout_reg[5] , 
        \tx_dout_reg[4] , \tx_dout_reg[3] , \tx_dout_reg[2] , 
        \tx_dout_reg[1] , \tx_dout_reg[0] }), .tx_hold_reg({
        \tx_hold_reg[7]_net_1 , \tx_hold_reg[6]_net_1 , 
        \tx_hold_reg[5]_net_1 , \tx_hold_reg[4]_net_1 , 
        \tx_hold_reg[3]_net_1 , \tx_hold_reg[2]_net_1 , 
        \tx_hold_reg[1]_net_1 , \tx_hold_reg[0]_net_1 }), 
        .fifo_write_tx(fifo_write_tx_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_full_tx_i_0(
        fifo_full_tx_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[3]  (.A(\rx_byte[3] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[3]_net_1 ), .Y(
        data_out[3]));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE clear_framing_error_reg0 (.D(clear_parity_en), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(clear_parity_reg0));
    SLE \tx_hold_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(GL0_INST), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[5]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_5), .Y(
        \rx_byte_in[5]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \genblk1.RXRDY5  (.A(rx_idle), .B(
        stop_strobe), .C(rx_dout_reg_empty_net_1), .Y(RXRDY5));
    CFG4 #( .INIT(16'h0004) )  fifo_read_rx_0_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(
        fifo_read_rx_0_sqmuxa));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[4]  (.A(\rx_byte[4] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[4]_net_1 ), .Y(
        data_out[4]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[2]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_2), .Y(
        \rx_byte_in[2]_net_1 ));
    mss_sb_CoreUARTapb_2_1_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s make_TX (
        .tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .counter({\counter[6] , \counter[5] , \counter[4] , 
        \counter[3] , \counter[2] , \counter[1] , \counter[0] }), 
        .controlReg2({controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .N_110(N_110)
        , .GPS_RX_c(GPS_RX_c), .CoreUARTapb_2_1_TXRDY(
        CoreUARTapb_2_1_TXRDY), .fifo_full_tx_i_0(fifo_full_tx_i_0), 
        .xmit_clock(xmit_clock), .baud_clock(baud_clock));
    SLE \tx_hold_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[6]_net_1 ));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[4]_net_1 ));
    mss_sb_CoreUARTapb_2_1_Clock_gen_0s make_CLOCK_GEN (.controlReg1({
        controlReg1[7], controlReg1[6], controlReg1[5], controlReg1[4], 
        controlReg1[3], controlReg1[2], controlReg1[1], controlReg1[0]})
        , .controlReg2({controlReg2[7], controlReg2[6], controlReg2[5], 
        controlReg2[4], controlReg2[3]}), .xmit_clock(xmit_clock), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .N_110(N_110));
    SLE \rx_state[1]  (.D(N_143_i), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_7));
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_1));
    CFG4 #( .INIT(16'hECCC) )  un1_clear_overflow (.A(un1_OEn_2), .B(
        overflow_reg5_net_1), .C(CoreAPB3_0_APBmslave3_PSELx), .D(
        un1_OEn_1), .Y(un1_clear_overflow_0));
    SLE clear_parity_reg (.D(clear_parity_reg0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_reg_net_1));
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_5));
    SLE overflow_reg (.D(overflow_reg5_net_1), .CLK(GL0_INST), .EN(
        un1_clear_overflow_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreUARTapb_2_1_OVERFLOW));
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_6));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \tx_hold_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[7]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(GL0_INST), 
        .EN(RXRDY5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_1_RXRDY));
    mss_sb_CoreUARTapb_2_1_fifo_256x8_0 \genblk3.rx_fifo  (.rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_byte_in({\rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte_in[4]_net_1 , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[1]_net_1 , \rx_byte_in[0]_net_1 }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_2318_i_0(N_2318_i_0), .N_2319_i_0(
        N_2319_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1_net_1), .fifo_full_rx(
        fifo_full_rx), .fifo_empty_rx(fifo_empty_rx));
    SLE \tx_hold_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[3]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \reg_write.tx_hold_reg5_i_0  (.A(un1_WEn_1)
        , .B(CoreAPB3_0_APBmslave3_PSELx), .C(un1_WEn_0), .Y(
        tx_hold_reg5_i_0));
    SLE fifo_write_tx (.D(tx_hold_reg5_i_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_write_tx_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[6]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_6), .Y(
        \rx_byte_in[6]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[7]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_7), .Y(
        \rx_byte_in[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[3]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[3] ), .Y(
        \rx_byte_in[3]_net_1 ));
    SLE \tx_hold_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hB333) )  rx_dout_reg_empty_1_sqmuxa_i (.A(
        un1_OEn_2), .B(rx_dout_reg4), .C(CoreAPB3_0_APBmslave3_PSELx), 
        .D(un1_OEn_1), .Y(rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_2));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[4]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[4] ), .Y(
        \rx_byte_in[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[0]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_0), .Y(
        \rx_byte_in[0]_net_1 ));
    SLE \tx_hold_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \reg_write.tx_hold_reg5  (.A(un1_WEn_1), 
        .B(CoreAPB3_0_APBmslave3_PSELx), .C(un1_WEn_0), .Y(
        tx_hold_reg5));
    
endmodule


module 
        mss_sb_CoreUARTapb_2_1_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s(
        
       CoreAPB3_0_APBmslave0_PWDATA,
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       un3_PRDATA_regif_1,
       CoreUARTapb_2_1_PARITY_ERR,
       N_97_1,
       CoreUARTapb_2_1_RXRDY,
       CoreUARTapb_2_1_TXRDY,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_0_APBmslave0_PENABLE,
       controlReg14_0,
       controlReg24_0,
       CoreAPB3_0_APBmslave0_PWRITE,
       psh_negedge_reg_1_sqmuxa_3_2,
       CoreUARTapb_2_1_FRAMING_ERR,
       CoreUARTapb_2_1_OVERFLOW,
       un1_WEn_1,
       un1_WEn_0,
       un1_OEn_2,
       un1_OEn_1,
       GPS_RX_c,
       GPS_TX_c
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [4:2] CoreAPB3_0_APBmslave0_PADDR;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  un3_PRDATA_regif_1;
output CoreUARTapb_2_1_PARITY_ERR;
input  N_97_1;
output CoreUARTapb_2_1_RXRDY;
output CoreUARTapb_2_1_TXRDY;
input  CoreAPB3_0_APBmslave3_PSELx;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  controlReg14_0;
input  controlReg24_0;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  psh_negedge_reg_1_sqmuxa_3_2;
output CoreUARTapb_2_1_FRAMING_ERR;
output CoreUARTapb_2_1_OVERFLOW;
input  un1_WEn_1;
input  un1_WEn_0;
input  un1_OEn_2;
input  un1_OEn_1;
output GPS_RX_c;
input  GPS_TX_c;

    wire \controlReg1[4]_net_1 , VCC_net_1, controlReg14, GND_net_1, 
        \controlReg1[5]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[7]_net_1 , \NxtPrdata[5] , un1_NxtPrdata23_i_0, 
        \NxtPrdata[6] , \NxtPrdata[7] , \controlReg2[0]_net_1 , 
        controlReg24, \controlReg2[1]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[7]_net_1 , \controlReg1[0]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[3]_net_1 , \NxtPrdata[0] , \NxtPrdata[1] , 
        \NxtPrdata[2] , \NxtPrdata[3] , \NxtPrdata[4] , 
        \NxtPrdata_5_bm[3]_net_1 , \NxtPrdata_5_am[3]_net_1 , 
        \NxtPrdata_5_bm[4]_net_1 , \NxtPrdata_5_am[4]_net_1 , 
        \NxtPrdata_5_bm[7]_net_1 , \NxtPrdata_5_am[7]_net_1 , 
        \NxtPrdata_5_bm[6]_net_1 , \NxtPrdata_5_am[6]_net_1 , 
        \NxtPrdata_5_bm[5]_net_1 , \NxtPrdata_5_am[5]_net_1 , N_275, 
        N_274, N_196, N_179, N_176, \rx_byte[0] , \rx_dout_reg[0] , 
        N_198, \rx_byte[2] , \rx_dout_reg[2] , N_181, \rx_byte[1] , 
        \rx_dout_reg[1] , N_178, \rx_dout_reg[5] , \rx_byte[5] , 
        \rx_dout_reg[6] , \rx_byte[6] , \rx_dout_reg[7] , \rx_byte[7] , 
        \data_out[4] , \data_out[3] ;
    
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[4]  (.A(
        CoreUARTapb_2_1_FRAMING_ERR), .B(\data_out[4] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[4]_net_1 ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[5]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[5] ), 
        .D(\rx_byte[5] ), .Y(\NxtPrdata_5_am[5]_net_1 ));
    SLE \controlReg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[5]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_1[2]  (.A(
        \rx_byte[2] ), .B(\rx_dout_reg[2] ), .C(N_274), .D(
        CoreUARTapb_2_1_PARITY_ERR), .Y(N_181));
    CFG4 #( .INIT(16'hFEEE) )  \NxtPrdata_5_0[0]  (.A(N_196), .B(N_198)
        , .C(CoreUARTapb_2_1_TXRDY), .D(N_275), .Y(\NxtPrdata[0] ));
    SLE \controlReg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[7]_net_1 ));
    SLE \iPRDATA[1]  (.D(\NxtPrdata[1] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[1]));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[6]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[6] ), 
        .D(\rx_byte[6] ), .Y(\NxtPrdata_5_am[6]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[7]  (.A(
        \controlReg2[7]_net_1 ), .B(\controlReg1[7]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[7]_net_1 ));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[1]  (.A(
        \controlReg1[1]_net_1 ), .B(\controlReg2[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_176));
    SLE \controlReg2[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[4]_net_1 ));
    SLE \iPRDATA[4]  (.D(\NxtPrdata[4] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[4]));
    VCC VCC (.Y(VCC_net_1));
    SLE \iPRDATA[3]  (.D(\NxtPrdata[3] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[3]));
    SLE \controlReg2[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[6]_net_1 ));
    SLE \controlReg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg1Seq.controlReg14  (.A(
        CoreAPB3_0_APBmslave3_PSELx), .B(CoreAPB3_0_APBmslave0_PENABLE)
        , .C(controlReg14_0), .Y(controlReg14));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[4]  (.A(
        \controlReg2[4]_net_1 ), .B(\controlReg1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[4]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[3]  (.A(
        CoreUARTapb_2_1_OVERFLOW), .B(\data_out[3] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[5]  (.A(
        \controlReg2[5]_net_1 ), .B(\controlReg1[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[5]_net_1 ));
    SLE \controlReg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[6]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_1[0]  (.A(
        \rx_byte[0] ), .B(\rx_dout_reg[0] ), .C(N_274), .D(
        CoreUARTapb_2_1_PARITY_ERR), .Y(N_198));
    SLE \controlReg2[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[3]_net_1 ));
    SLE \controlReg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[2]_net_1 ));
    SLE \controlReg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[4]_net_1 ));
    SLE \iPRDATA[5]  (.D(\NxtPrdata[5] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[5]));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[0]  (.A(
        \controlReg1[0]_net_1 ), .B(\controlReg2[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_196));
    SLE \iPRDATA[7]  (.D(\NxtPrdata[7] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[7]));
    SLE \controlReg2[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[1]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[6]  (.A(
        \controlReg2[6]_net_1 ), .B(\controlReg1[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[6]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[4]_net_1 ), 
        .C(\NxtPrdata_5_am[4]_net_1 ), .Y(\NxtPrdata[4] ));
    SLE \controlReg2[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[7]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24  (.A(
        CoreAPB3_0_APBmslave3_PSELx), .B(CoreAPB3_0_APBmslave0_PENABLE)
        , .C(controlReg24_0), .Y(controlReg24));
    SLE \iPRDATA[2]  (.D(\NxtPrdata[2] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[2]));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[3]_net_1 ), 
        .C(\NxtPrdata_5_am[3]_net_1 ), .Y(\NxtPrdata[3] ));
    SLE \controlReg2[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[5]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[3]  (.A(
        \controlReg2[3]_net_1 ), .B(\controlReg1[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[3]_net_1 ));
    SLE \controlReg2[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[2]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  un1_NxtPrdata23_i (.A(
        CoreAPB3_0_APBmslave0_PWRITE), .B(
        CoreAPB3_0_APBmslave0_PENABLE), .C(
        psh_negedge_reg_1_sqmuxa_3_2), .D(CoreAPB3_0_APBmslave3_PSELx), 
        .Y(un1_NxtPrdata23_i_0));
    SLE \iPRDATA[6]  (.D(\NxtPrdata[6] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[6]));
    SLE \iPRDATA[0]  (.D(\NxtPrdata[0] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreAPB3_0_APBmslave3_PRDATA[0]));
    mss_sb_CoreUARTapb_2_1_COREUART_1s_1s_0s_15s_0s uUART (
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .data_out({\data_out[4] , 
        \data_out[3] }), .controlReg1({\controlReg1[7]_net_1 , 
        \controlReg1[6]_net_1 , \controlReg1[5]_net_1 , 
        \controlReg1[4]_net_1 , \controlReg1[3]_net_1 , 
        \controlReg1[2]_net_1 , \controlReg1[1]_net_1 , 
        \controlReg1[0]_net_1 }), .controlReg2({\controlReg2[7]_net_1 , 
        \controlReg2[6]_net_1 , \controlReg2[5]_net_1 , 
        \controlReg2[4]_net_1 , \controlReg2[3]_net_1 , 
        \controlReg2[2]_net_1 , \controlReg2[1]_net_1 , 
        \controlReg2[0]_net_1 }), .rx_dout_reg_5(\rx_dout_reg[5] ), 
        .rx_dout_reg_6(\rx_dout_reg[6] ), .rx_dout_reg_7(
        \rx_dout_reg[7] ), .rx_dout_reg_0(\rx_dout_reg[0] ), 
        .rx_dout_reg_1(\rx_dout_reg[1] ), .rx_dout_reg_2(
        \rx_dout_reg[2] ), .rx_byte_5(\rx_byte[5] ), .rx_byte_0(
        \rx_byte[0] ), .rx_byte_2(\rx_byte[2] ), .rx_byte_1(
        \rx_byte[1] ), .rx_byte_6(\rx_byte[6] ), .rx_byte_7(
        \rx_byte[7] ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreUARTapb_2_1_OVERFLOW(CoreUARTapb_2_1_OVERFLOW), 
        .CoreUARTapb_2_1_RXRDY(CoreUARTapb_2_1_RXRDY), .un1_WEn_1(
        un1_WEn_1), .CoreAPB3_0_APBmslave3_PSELx(
        CoreAPB3_0_APBmslave3_PSELx), .un1_WEn_0(un1_WEn_0), 
        .CoreUARTapb_2_1_PARITY_ERR(CoreUARTapb_2_1_PARITY_ERR), 
        .un1_OEn_2(un1_OEn_2), .un1_OEn_1(un1_OEn_1), .GPS_RX_c(
        GPS_RX_c), .CoreUARTapb_2_1_TXRDY(CoreUARTapb_2_1_TXRDY), 
        .GPS_TX_c(GPS_TX_c), .CoreUARTapb_2_1_FRAMING_ERR(
        CoreUARTapb_2_1_FRAMING_ERR));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[7]_net_1 ), 
        .C(\NxtPrdata_5_am[7]_net_1 ), .Y(\NxtPrdata[7] ));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[2]  (.A(
        \controlReg1[2]_net_1 ), .B(\controlReg2[2]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_179));
    CFG2 #( .INIT(4'h4) )  \NxtPrdata_5_0_a2_2[1]  (.A(
        un3_PRDATA_regif_1), .B(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        N_274));
    CFG4 #( .INIT(16'hFEEE) )  \NxtPrdata_5_0[2]  (.A(N_179), .B(N_181)
        , .C(CoreUARTapb_2_1_PARITY_ERR), .D(N_275), .Y(\NxtPrdata[2] )
        );
    SLE \controlReg2[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[0]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[6]_net_1 ), 
        .C(\NxtPrdata_5_am[6]_net_1 ), .Y(\NxtPrdata[6] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[7]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_97_1), .C(\rx_dout_reg[7] ), 
        .D(\rx_byte[7] ), .Y(\NxtPrdata_5_am[7]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_1[1]  (.A(
        \rx_byte[1] ), .B(\rx_dout_reg[1] ), .C(N_274), .D(
        CoreUARTapb_2_1_PARITY_ERR), .Y(N_178));
    CFG3 #( .INIT(8'h04) )  \NxtPrdata_5_0_a2_3[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_275));
    SLE \controlReg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[1]_net_1 ));
    CFG4 #( .INIT(16'hFEEE) )  \NxtPrdata_5_0[1]  (.A(N_176), .B(N_178)
        , .C(CoreUARTapb_2_1_RXRDY), .D(N_275), .Y(\NxtPrdata[1] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[5]_net_1 ), 
        .C(\NxtPrdata_5_am[5]_net_1 ), .Y(\NxtPrdata[5] ));
    SLE \controlReg1[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[0]_net_1 ));
    
endmodule


module pwm_gen_10s_16s_0(
       PWM_c,
       period_cnt,
       pwm_negedge_reg,
       pwm_enable_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST
    );
output [10:1] PWM_c;
input  [15:0] period_cnt;
input  [160:1] pwm_negedge_reg;
input  [10:1] pwm_enable_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;

    wire VCC_net_1, \PWM_int_38[3] , \un1_pwm_enable_reg_9_i_0[0] , 
        GND_net_1, \PWM_int_24[2] , \un1_pwm_enable_reg_6_i_0[0] , 
        \PWM_int_10[1] , \un1_pwm_enable_reg_7_i_0[0] , 
        \PWM_int_136[10] , \un1_pwm_enable_reg_i_0[0] , 
        \PWM_int_122[9] , \un1_pwm_enable_reg_1_i_0[0] , 
        \PWM_int_108[8] , \un1_pwm_enable_reg_4_i_0[0] , N_29_i_0, N_5, 
        \PWM_int_80[6] , \un1_pwm_enable_reg_2_i_0[0] , N_31_i_0, N_7, 
        \PWM_int_52[4] , \un1_pwm_enable_reg_8_i_0[0] , 
        \un1_period_cnt_1_1_data_tmp[0] , 
        \un1_period_cnt_1_1_data_tmp[1] , 
        \un1_period_cnt_1_1_data_tmp[2] , 
        \un1_period_cnt_1_1_data_tmp[3] , 
        \un1_period_cnt_1_1_data_tmp[4] , 
        \un1_period_cnt_1_1_data_tmp[5] , 
        \un1_period_cnt_1_1_data_tmp[6] , un1_period_cnt_1, 
        \un1_period_cnt_1_0_data_tmp[0] , 
        \un1_period_cnt_1_0_data_tmp[1] , 
        \un1_period_cnt_1_0_data_tmp[2] , 
        \un1_period_cnt_1_0_data_tmp[3] , 
        \un1_period_cnt_1_0_data_tmp[4] , 
        \un1_period_cnt_1_0_data_tmp[5] , 
        \un1_period_cnt_1_0_data_tmp[6] , un1_period_cnt_1_0, 
        \un1_period_cnt_1_0_data_tmp_0[0] , 
        \un1_period_cnt_1_0_data_tmp_0[1] , 
        \un1_period_cnt_1_0_data_tmp_0[2] , 
        \un1_period_cnt_1_0_data_tmp_0[3] , 
        \un1_period_cnt_1_0_data_tmp_0[4] , 
        \un1_period_cnt_1_0_data_tmp_0[5] , 
        \un1_period_cnt_1_0_data_tmp_0[6] , un1_period_cnt_1_1, 
        \un1_period_cnt_1_0_data_tmp_1[0] , 
        \un1_period_cnt_1_0_data_tmp_1[1] , 
        \un1_period_cnt_1_0_data_tmp_1[2] , 
        \un1_period_cnt_1_0_data_tmp_1[3] , 
        \un1_period_cnt_1_0_data_tmp_1[4] , 
        \un1_period_cnt_1_0_data_tmp_1[5] , 
        \un1_period_cnt_1_0_data_tmp_1[6] , un1_period_cnt_1_2, 
        \un1_period_cnt_1_0_data_tmp_2[0] , 
        \un1_period_cnt_1_0_data_tmp_2[1] , 
        \un1_period_cnt_1_0_data_tmp_2[2] , 
        \un1_period_cnt_1_0_data_tmp_2[3] , 
        \un1_period_cnt_1_0_data_tmp_2[4] , 
        \un1_period_cnt_1_0_data_tmp_2[5] , 
        \un1_period_cnt_1_0_data_tmp_2[6] , un1_period_cnt_1_3, 
        \un1_period_cnt_1_0_data_tmp_3[0] , 
        \un1_period_cnt_1_0_data_tmp_3[1] , 
        \un1_period_cnt_1_0_data_tmp_3[2] , 
        \un1_period_cnt_1_0_data_tmp_3[3] , 
        \un1_period_cnt_1_0_data_tmp_3[4] , 
        \un1_period_cnt_1_0_data_tmp_3[5] , 
        \un1_period_cnt_1_0_data_tmp_3[6] , un1_period_cnt_1_4, 
        \un1_period_cnt_1_0_data_tmp_4[0] , 
        \un1_period_cnt_1_0_data_tmp_4[1] , 
        \un1_period_cnt_1_0_data_tmp_4[2] , 
        \un1_period_cnt_1_0_data_tmp_4[3] , 
        \un1_period_cnt_1_0_data_tmp_4[4] , 
        \un1_period_cnt_1_0_data_tmp_4[5] , 
        \un1_period_cnt_1_0_data_tmp_4[6] , un1_period_cnt_1_5, 
        \un1_period_cnt_1_0_data_tmp_5[0] , 
        \un1_period_cnt_1_0_data_tmp_5[1] , 
        \un1_period_cnt_1_0_data_tmp_5[2] , 
        \un1_period_cnt_1_0_data_tmp_5[3] , 
        \un1_period_cnt_1_0_data_tmp_5[4] , 
        \un1_period_cnt_1_0_data_tmp_5[5] , 
        \un1_period_cnt_1_0_data_tmp_5[6] , un1_period_cnt_1_6, 
        \un1_period_cnt_1_0_data_tmp_6[0] , 
        \un1_period_cnt_1_0_data_tmp_6[1] , 
        \un1_period_cnt_1_0_data_tmp_6[2] , 
        \un1_period_cnt_1_0_data_tmp_6[3] , 
        \un1_period_cnt_1_0_data_tmp_6[4] , 
        \un1_period_cnt_1_0_data_tmp_6[5] , 
        \un1_period_cnt_1_0_data_tmp_6[6] , un1_period_cnt_1_7, 
        \un1_period_cnt_1_0_data_tmp_7[0] , 
        \un1_period_cnt_1_0_data_tmp_7[1] , 
        \un1_period_cnt_1_0_data_tmp_7[2] , 
        \un1_period_cnt_1_0_data_tmp_7[3] , 
        \un1_period_cnt_1_0_data_tmp_7[4] , 
        \un1_period_cnt_1_0_data_tmp_7[5] , 
        \un1_period_cnt_1_0_data_tmp_7[6] , un1_period_cnt_1_8, 
        \PWM_int_24_f1_2[2] , \PWM_int_136_f1_2[10] , 
        \PWM_int_80_f1_2[6] , \PWM_int_52_f1_2[4] , 
        \PWM_int_108_f1_2[8] , \PWM_int_10_f1_2[1] , 
        \PWM_int_122_f1_2[9] , \PWM_int_38_f1_2[3] , 
        \PWM_int_66_f0_i_3_3[5] , \PWM_int_24_f1_11[2] , 
        \PWM_int_24_f1_10[2] , \PWM_int_24_f1_8[2] , 
        \PWM_int_136_f1_11[10] , \PWM_int_136_f1_10[10] , 
        \PWM_int_136_f1_8[10] , \PWM_int_80_f1_11[6] , 
        \PWM_int_80_f1_10[6] , \PWM_int_80_f1_8[6] , 
        \PWM_int_52_f1_11[4] , \PWM_int_52_f1_10[4] , 
        \PWM_int_52_f1_8[4] , \PWM_int_108_f1_11[8] , 
        \PWM_int_108_f1_10[8] , \PWM_int_108_f1_8[8] , 
        \PWM_int_10_f1_11[1] , \PWM_int_10_f1_10[1] , 
        \PWM_int_10_f1_8[1] , \PWM_int_122_f1_11[9] , 
        \PWM_int_122_f1_10[9] , \PWM_int_122_f1_8[9] , 
        \PWM_int_66_f0_i_a9_11[5] , \PWM_int_66_f0_i_a9_10[5] , 
        \PWM_int_66_f0_i_a9_9[5] , \PWM_int_66_f0_i_a9_8[5] , 
        \PWM_int_38_f1_11[3] , \PWM_int_38_f1_10[3] , 
        \PWM_int_38_f1_8[3] , \PWM_int_94_f0_i_a9_11[7] , 
        \PWM_int_94_f0_i_a9_10[7] , \PWM_int_94_f0_i_a9_9[7] , 
        \PWM_int_94_f0_i_a9_8[7] , \PWM_int_66_f0_i_3_4[5] , N_29_1, 
        N_29_2, \PWM_int_24_f1_13[2] , \PWM_int_136_f1_13[10] , 
        \PWM_int_80_f1_13[6] , \PWM_int_52_f1_13[4] , 
        \PWM_int_108_f1_13[8] , \PWM_int_10_f1_13[1] , 
        \PWM_int_122_f1_13[9] , \PWM_int_38_f1_13[3] , N_29_3, 
        \PWM_int_24_f1_14[2] , \PWM_int_136_f1_14[10] , 
        \PWM_int_80_f1_14[6] , \PWM_int_52_f1_14[4] , 
        \PWM_int_108_f1_14[8] , \PWM_int_10_f1_14[1] , 
        \PWM_int_122_f1_14[9] , \PWM_int_66_f0_i_a9_14[5] , 
        \PWM_int_38_f1_14[3] , \PWM_int_94_f0_i_a9_14[7] , 
        un1_period_cnt_NE_i_0, \PWM_int_94_f0_i_1[7] , 
        \PWM_int_66_f0_i_1[5] ;
    
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[42]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[41]), .FCI(\un1_period_cnt_1_0_data_tmp_7[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_7[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_14[6]  (.A(
        pwm_negedge_reg[83]), .B(pwm_negedge_reg[82]), .C(
        \PWM_int_80_f1_11[6] ), .D(\PWM_int_80_f1_8[6] ), .Y(
        \PWM_int_80_f1_14[6] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_14[3]  (.A(
        pwm_negedge_reg[35]), .B(pwm_negedge_reg[34]), .C(
        \PWM_int_38_f1_11[3] ), .D(\PWM_int_38_f1_8[3] ), .Y(
        \PWM_int_38_f1_14[3] ));
    SLE \PWM_output_generation[1].genblk1.PWM_int[1]  (.D(
        \PWM_int_10[1] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_7_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[1]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[140]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[139]), .FCI(
        \un1_period_cnt_1_0_data_tmp[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[5] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a9_14[7]  (
        .A(pwm_negedge_reg[101]), .B(pwm_negedge_reg[98]), .C(
        \PWM_int_94_f0_i_a9_11[7] ), .D(\PWM_int_94_f0_i_a9_8[7] ), .Y(
        \PWM_int_94_f0_i_a9_14[7] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[120]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[119]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_10[4]  (.A(
        pwm_negedge_reg[64]), .B(pwm_negedge_reg[59]), .C(
        pwm_negedge_reg[57]), .D(pwm_negedge_reg[56]), .Y(
        \PWM_int_52_f1_10[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_14[8]  (.A(
        pwm_negedge_reg[118]), .B(pwm_negedge_reg[116]), .C(
        \PWM_int_108_f1_11[8] ), .D(\PWM_int_108_f1_8[8] ), .Y(
        \PWM_int_108_f1_14[8] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_11[10]  (.A(
        pwm_negedge_reg[151]), .B(pwm_negedge_reg[150]), .C(
        pwm_negedge_reg[149]), .D(pwm_negedge_reg[148]), .Y(
        \PWM_int_136_f1_11[10] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f0[4]  (.A(
        \PWM_int_52_f1_14[4] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[4]), .D(\PWM_int_52_f1_13[4] ), .Y(
        \PWM_int_52[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[40]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[39]), .FCI(\un1_period_cnt_1_0_data_tmp_7[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_7[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[102]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[101]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[98]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[97]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_1[5]  (.A(
        period_cnt[5]), .B(period_cnt[4]), .C(period_cnt[3]), .D(
        period_cnt[2]), .Y(N_29_1));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_2[6]  (.A(
        pwm_negedge_reg[92]), .B(pwm_negedge_reg[93]), .Y(
        \PWM_int_80_f1_2[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[108]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[107]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[5] ));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a9_8[7]  (.A(
        pwm_negedge_reg[103]), .B(pwm_negedge_reg[97]), .C(PWM_c[7]), 
        .Y(\PWM_int_94_f0_i_a9_8[7] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_13[10]  (.A(
        pwm_negedge_reg[152]), .B(pwm_negedge_reg[153]), .C(
        \PWM_int_136_f1_10[10] ), .D(\PWM_int_136_f1_2[10] ), .Y(
        \PWM_int_136_f1_13[10] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_11[1]  (.A(
        pwm_negedge_reg[4]), .B(pwm_negedge_reg[3]), .C(
        pwm_negedge_reg[2]), .D(pwm_negedge_reg[1]), .Y(
        \PWM_int_10_f1_11[1] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[8].genblk1.PWM_int_RNO[8]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[8]), .C(
        un1_period_cnt_1_5), .Y(\un1_pwm_enable_reg_4_i_0[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_15  (
        .A(pwm_negedge_reg[156]), .B(period_cnt[10]), .C(
        period_cnt[11]), .D(pwm_negedge_reg[155]), .FCI(
        \un1_period_cnt_1_1_data_tmp[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_9  (.A(
        pwm_negedge_reg[158]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[157]), .FCI(
        \un1_period_cnt_1_1_data_tmp[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[6] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_11[6]  (.A(
        pwm_negedge_reg[87]), .B(pwm_negedge_reg[86]), .C(
        pwm_negedge_reg[85]), .D(pwm_negedge_reg[84]), .Y(
        \PWM_int_80_f1_11[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[62]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[61]), .FCI(
        \un1_period_cnt_1_0_data_tmp_6[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_6[6] ));
    SLE \PWM_output_generation[3].genblk1.PWM_int[3]  (.D(
        \PWM_int_38[3] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_9_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[3]));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_2[9]  (.A(
        pwm_negedge_reg[129]), .B(pwm_negedge_reg[132]), .Y(
        \PWM_int_122_f1_2[9] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_2[4]  (.A(
        pwm_negedge_reg[58]), .B(pwm_negedge_reg[61]), .Y(
        \PWM_int_52_f1_2[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_10[10]  (.A(
        pwm_negedge_reg[159]), .B(pwm_negedge_reg[158]), .C(
        pwm_negedge_reg[157]), .D(pwm_negedge_reg[156]), .Y(
        \PWM_int_136_f1_10[10] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[3].genblk1.PWM_int_RNO[3]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[3]), .C(
        un1_period_cnt_1_8), .Y(\un1_pwm_enable_reg_9_i_0[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_13[4]  (.A(
        pwm_negedge_reg[60]), .B(pwm_negedge_reg[63]), .C(
        \PWM_int_52_f1_10[4] ), .D(\PWM_int_52_f1_2[4] ), .Y(
        \PWM_int_52_f1_13[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[10]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[9]), .FCI(\un1_period_cnt_1_0_data_tmp_1[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[4] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_8[8]  (.A(
        pwm_negedge_reg[127]), .B(pwm_negedge_reg[117]), .C(PWM_c[8]), 
        .Y(\PWM_int_108_f1_8[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[16]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[15]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_2));
    SLE \PWM_output_generation[10].genblk1.PWM_int[10]  (.D(
        \PWM_int_136[10] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_i_0[0] ), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[10]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_14[2]  (.A(
        pwm_negedge_reg[22]), .B(pwm_negedge_reg[21]), .C(
        \PWM_int_24_f1_11[2] ), .D(\PWM_int_24_f1_8[2] ), .Y(
        \PWM_int_24_f1_14[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_27  (
        .A(pwm_negedge_reg[154]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[153]), .FCI(
        \un1_period_cnt_1_1_data_tmp[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_13[9]  (.A(
        pwm_negedge_reg[130]), .B(pwm_negedge_reg[131]), .C(
        \PWM_int_122_f1_10[9] ), .D(\PWM_int_122_f1_2[9] ), .Y(
        \PWM_int_122_f1_13[9] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_2[3]  (.A(
        pwm_negedge_reg[41]), .B(pwm_negedge_reg[47]), .Y(
        \PWM_int_38_f1_2[3] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0[2]  (.A(
        \PWM_int_24_f1_14[2] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[2]), .D(\PWM_int_24_f1_13[2] ), .Y(
        \PWM_int_24[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[50]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[49]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_6[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[132]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[131]), .FCI(
        \un1_period_cnt_1_0_data_tmp[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[52]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[51]), .FCI(\un1_period_cnt_1_0_data_tmp_6[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_6[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[32]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[31]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_1));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f0[10]  (.A(
        \PWM_int_136_f1_14[10] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[10]), .D(\PWM_int_136_f1_13[10] ), .Y(
        \PWM_int_136[10] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_13[8]  (.A(
        pwm_negedge_reg[124]), .B(pwm_negedge_reg[126]), .C(
        \PWM_int_108_f1_10[8] ), .D(\PWM_int_108_f1_2[8] ), .Y(
        \PWM_int_108_f1_13[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[8]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[7]), .FCI(\un1_period_cnt_1_0_data_tmp_1[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[106]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[105]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_11[9]  (.A(
        pwm_negedge_reg[139]), .B(pwm_negedge_reg[138]), .C(
        pwm_negedge_reg[137]), .D(pwm_negedge_reg[136]), .Y(
        \PWM_int_122_f1_11[9] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[60]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[59]), .FCI(
        \un1_period_cnt_1_0_data_tmp_6[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_6[5] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[2].genblk1.PWM_int_RNO[2]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[2]), .C(
        un1_period_cnt_1_1), .Y(\un1_pwm_enable_reg_6_i_0[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[116]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[115]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_10[2]  (.A(
        pwm_negedge_reg[32]), .B(pwm_negedge_reg[31]), .C(
        pwm_negedge_reg[30]), .D(pwm_negedge_reg[29]), .Y(
        \PWM_int_24_f1_10[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_11[3]  (.A(
        pwm_negedge_reg[39]), .B(pwm_negedge_reg[38]), .C(
        pwm_negedge_reg[37]), .D(pwm_negedge_reg[36]), .Y(
        \PWM_int_38_f1_11[3] ));
    CFG3 #( .INIT(8'hFB) )  \un1_pwm_enable_reg_5_i_0[0]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[7]), .C(
        un1_period_cnt_1_6), .Y(N_5));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[104]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[103]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_2[5]  (.A(
        period_cnt[7]), .B(period_cnt[6]), .C(period_cnt[1]), .D(
        period_cnt[0]), .Y(N_29_2));
    SLE \PWM_output_generation[2].genblk1.PWM_int[2]  (.D(
        \PWM_int_24[2] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_6_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[2]));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_13[3]  (.A(
        pwm_negedge_reg[40]), .B(pwm_negedge_reg[43]), .C(
        \PWM_int_38_f1_10[3] ), .D(\PWM_int_38_f1_2[3] ), .Y(
        \PWM_int_38_f1_13[3] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_8[9]  (.A(
        pwm_negedge_reg[143]), .B(pwm_negedge_reg[142]), .C(PWM_c[9]), 
        .Y(\PWM_int_122_f1_8[9] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[46]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[45]), .FCI(
        \un1_period_cnt_1_0_data_tmp_7[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_7[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[84]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[83]), .FCI(\un1_period_cnt_1_0_data_tmp_2[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_11[8]  (.A(
        pwm_negedge_reg[119]), .B(pwm_negedge_reg[115]), .C(
        pwm_negedge_reg[114]), .D(pwm_negedge_reg[113]), .Y(
        \PWM_int_108_f1_11[8] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_14[9]  (.A(
        pwm_negedge_reg[141]), .B(pwm_negedge_reg[140]), .C(
        \PWM_int_122_f1_11[9] ), .D(\PWM_int_122_f1_8[9] ), .Y(
        \PWM_int_122_f1_14[9] ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_a9_8[5]  (.A(
        pwm_negedge_reg[79]), .B(pwm_negedge_reg[78]), .C(PWM_c[5]), 
        .Y(\PWM_int_66_f0_i_a9_8[5] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_11[4]  (.A(
        pwm_negedge_reg[55]), .B(pwm_negedge_reg[51]), .C(
        pwm_negedge_reg[50]), .D(pwm_negedge_reg[49]), .Y(
        \PWM_int_52_f1_11[4] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_2[10]  (.A(
        pwm_negedge_reg[154]), .B(pwm_negedge_reg[155]), .Y(
        \PWM_int_136_f1_2[10] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_10[1]  (.A(
        pwm_negedge_reg[12]), .B(pwm_negedge_reg[11]), .C(
        pwm_negedge_reg[10]), .D(pwm_negedge_reg[9]), .Y(
        \PWM_int_10_f1_10[1] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_a9_14[5]  (
        .A(pwm_negedge_reg[77]), .B(pwm_negedge_reg[76]), .C(
        \PWM_int_66_f0_i_a9_11[5] ), .D(\PWM_int_66_f0_i_a9_8[5] ), .Y(
        \PWM_int_66_f0_i_a9_14[5] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_a9_10[5]  (
        .A(pwm_negedge_reg[71]), .B(pwm_negedge_reg[70]), .C(
        pwm_negedge_reg[69]), .D(pwm_negedge_reg[68]), .Y(
        \PWM_int_66_f0_i_a9_10[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[90]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[89]), .FCI(\un1_period_cnt_1_0_data_tmp_2[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[36]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[35]), .FCI(\un1_period_cnt_1_0_data_tmp_7[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_7[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[142]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[141]), .FCI(
        \un1_period_cnt_1_0_data_tmp[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[6] ));
    SLE \PWM_output_generation[7].genblk1.PWM_int[7]  (.D(N_29_i_0), 
        .CLK(GL0_INST), .EN(N_5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[7]));
    SLE \PWM_output_generation[6].genblk1.PWM_int[6]  (.D(
        \PWM_int_80[6] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_2_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[6]));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_2[8]  (.A(
        pwm_negedge_reg[123]), .B(pwm_negedge_reg[125]), .Y(
        \PWM_int_108_f1_2[8] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_8[10]  (.A(
        pwm_negedge_reg[160]), .B(pwm_negedge_reg[145]), .C(PWM_c[10]), 
        .Y(\PWM_int_136_f1_8[10] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[134]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[133]), .FCI(
        \un1_period_cnt_1_0_data_tmp[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[88]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[87]), .FCI(\un1_period_cnt_1_0_data_tmp_2[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[3] ));
    SLE \PWM_output_generation[9].genblk1.PWM_int[9]  (.D(
        \PWM_int_122[9] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_1_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[9]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[112]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[111]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_6));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f0[6]  (.A(
        \PWM_int_80_f1_14[6] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[6]), .D(\PWM_int_80_f1_13[6] ), .Y(
        \PWM_int_80[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[54]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[53]), .FCI(\un1_period_cnt_1_0_data_tmp_6[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_6[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[34]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[33]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_7[0] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0[1]  (.A(
        \PWM_int_10_f1_14[1] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[1]), .D(\PWM_int_10_f1_13[1] ), .Y(
        \PWM_int_10[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[18]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[17]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_13[6]  (.A(
        pwm_negedge_reg[94]), .B(pwm_negedge_reg[95]), .C(
        \PWM_int_80_f1_10[6] ), .D(\PWM_int_80_f1_2[6] ), .Y(
        \PWM_int_80_f1_13[6] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_8[4]  (.A(
        pwm_negedge_reg[62]), .B(pwm_negedge_reg[53]), .C(PWM_c[4]), 
        .Y(\PWM_int_52_f1_8[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[118]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[117]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[44]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[43]), .FCI(
        \un1_period_cnt_1_0_data_tmp_7[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_7[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[20]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[19]), .FCI(\un1_period_cnt_1_0_data_tmp_0[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_0[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_11[2]  (.A(
        pwm_negedge_reg[20]), .B(pwm_negedge_reg[19]), .C(
        pwm_negedge_reg[18]), .D(pwm_negedge_reg[17]), .Y(
        \PWM_int_24_f1_11[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_14[1]  (.A(
        pwm_negedge_reg[6]), .B(pwm_negedge_reg[5]), .C(
        \PWM_int_10_f1_11[1] ), .D(\PWM_int_10_f1_8[1] ), .Y(
        \PWM_int_10_f1_14[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[28]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[27]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[14]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[13]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[86]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[85]), .FCI(\un1_period_cnt_1_0_data_tmp_2[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[66]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[65]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[110]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[109]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_1  (.A(
        pwm_negedge_reg[146]), .B(period_cnt[0]), .C(period_cnt[1]), 
        .D(pwm_negedge_reg[145]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[0] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[1].genblk1.PWM_int_RNO[1]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[1]), .C(
        un1_period_cnt_1_2), .Y(\un1_pwm_enable_reg_7_i_0[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[96]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[95]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_3));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[68]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[67]), .FCI(\un1_period_cnt_1_0_data_tmp_3[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[4]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[3]), .FCI(\un1_period_cnt_1_0_data_tmp_1[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[76]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[75]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[5] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_8[6]  (.A(
        pwm_negedge_reg[96]), .B(pwm_negedge_reg[81]), .C(PWM_c[6]), 
        .Y(\PWM_int_80_f1_8[6] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_2[1]  (.A(
        pwm_negedge_reg[13]), .B(pwm_negedge_reg[14]), .Y(
        \PWM_int_10_f1_2[1] ));
    SLE \PWM_output_generation[5].genblk1.PWM_int[5]  (.D(N_31_i_0), 
        .CLK(GL0_INST), .EN(N_7), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[5]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[38]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[37]), .FCI(\un1_period_cnt_1_0_data_tmp_7[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_7[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_33  (
        .A(pwm_negedge_reg[150]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[149]), .FCI(
        \un1_period_cnt_1_1_data_tmp[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_14[4]  (.A(
        pwm_negedge_reg[54]), .B(pwm_negedge_reg[52]), .C(
        \PWM_int_52_f1_11[4] ), .D(\PWM_int_52_f1_8[4] ), .Y(
        \PWM_int_52_f1_14[4] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f0[9]  (.A(
        \PWM_int_122_f1_14[9] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[9]), .D(\PWM_int_122_f1_13[9] ), .Y(
        \PWM_int_122[9] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a9_9[7]  (.A(
        pwm_negedge_reg[110]), .B(pwm_negedge_reg[109]), .C(
        pwm_negedge_reg[108]), .D(pwm_negedge_reg[102]), .Y(
        \PWM_int_94_f0_i_a9_9[7] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_45  (
        .A(pwm_negedge_reg[160]), .B(period_cnt[14]), .C(
        period_cnt[15]), .D(pwm_negedge_reg[159]), .FCI(
        \un1_period_cnt_1_1_data_tmp[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_8[2]  (.A(
        pwm_negedge_reg[24]), .B(pwm_negedge_reg[23]), .C(PWM_c[2]), 
        .Y(\PWM_int_24_f1_8[2] ));
    CFG4 #( .INIT(16'h1333) )  
        \PWM_output_generation[5].genblk1.PWM_int_RNO[5]  (.A(
        \PWM_int_66_f0_i_a9_14[5] ), .B(\PWM_int_66_f0_i_1[5] ), .C(
        \PWM_int_66_f0_i_a9_10[5] ), .D(\PWM_int_66_f0_i_a9_9[5] ), .Y(
        N_31_i_0));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[114]), .B(period_cnt[0]), .C(period_cnt[1]), 
        .D(pwm_negedge_reg[113]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[0] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_a9_11[5]  (
        .A(pwm_negedge_reg[75]), .B(pwm_negedge_reg[74]), .C(
        pwm_negedge_reg[73]), .D(pwm_negedge_reg[72]), .Y(
        \PWM_int_66_f0_i_a9_11[5] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a9_10[7]  (
        .A(pwm_negedge_reg[107]), .B(pwm_negedge_reg[106]), .C(
        pwm_negedge_reg[105]), .D(pwm_negedge_reg[104]), .Y(
        \PWM_int_94_f0_i_a9_10[7] ));
    CFG4 #( .INIT(16'hFFFB) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_1[7]  (.A(
        N_29_2), .B(pwm_enable_reg[7]), .C(N_29_3), .D(N_29_1), .Y(
        \PWM_int_94_f0_i_1[7] ));
    CFG3 #( .INIT(8'h01) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_1_RNIQ0711[5]  
        (.A(N_29_1), .B(N_29_3), .C(N_29_2), .Y(un1_period_cnt_NE_i_0));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[10].genblk1.PWM_int_136_f1_14[10]  (.A(
        pwm_negedge_reg[147]), .B(pwm_negedge_reg[146]), .C(
        \PWM_int_136_f1_11[10] ), .D(\PWM_int_136_f1_8[10] ), .Y(
        \PWM_int_136_f1_14[10] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[124]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[123]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[48]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[47]), .FCI(
        \un1_period_cnt_1_0_data_tmp_7[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_8));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[30]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[29]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[128]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[127]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_5));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_10[6]  (.A(
        pwm_negedge_reg[91]), .B(pwm_negedge_reg[90]), .C(
        pwm_negedge_reg[89]), .D(pwm_negedge_reg[88]), .Y(
        \PWM_int_80_f1_10[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[82]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[81]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[0] ));
    CFG4 #( .INIT(16'hFFFB) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_1_2[5]  (.A(
        N_29_2), .B(pwm_enable_reg[5]), .C(N_29_3), .D(N_29_1), .Y(
        \PWM_int_66_f0_i_1[5] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[9].genblk1.PWM_int_122_f1_10[9]  (.A(
        pwm_negedge_reg[144]), .B(pwm_negedge_reg[135]), .C(
        pwm_negedge_reg[134]), .D(pwm_negedge_reg[133]), .Y(
        \PWM_int_122_f1_10[9] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[22]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[21]), .FCI(\un1_period_cnt_1_0_data_tmp_0[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_0[2] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_a9_9[5]  (.A(
        pwm_negedge_reg[80]), .B(pwm_negedge_reg[67]), .C(
        pwm_negedge_reg[66]), .D(pwm_negedge_reg[65]), .Y(
        \PWM_int_66_f0_i_a9_9[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[74]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[73]), .FCI(\un1_period_cnt_1_0_data_tmp_3[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[4] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_3_3[5]  (.A(
        period_cnt[12]), .B(period_cnt[13]), .Y(
        \PWM_int_66_f0_i_3_3[5] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_13[2]  (.A(
        pwm_negedge_reg[25]), .B(pwm_negedge_reg[26]), .C(
        \PWM_int_24_f1_10[2] ), .D(\PWM_int_24_f1_2[2] ), .Y(
        \PWM_int_24_f1_13[2] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a9_11[7]  (
        .A(pwm_negedge_reg[112]), .B(pwm_negedge_reg[111]), .C(
        pwm_negedge_reg[100]), .D(pwm_negedge_reg[99]), .Y(
        \PWM_int_94_f0_i_a9_11[7] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[92]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[91]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[5] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[10].genblk1.PWM_int_RNO[10]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[10]), .C(
        un1_period_cnt_1), .Y(\un1_pwm_enable_reg_i_0[0] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_8[1]  (.A(
        pwm_negedge_reg[8]), .B(pwm_negedge_reg[7]), .C(PWM_c[1]), .Y(
        \PWM_int_10_f1_8[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[144]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[143]), .FCI(
        \un1_period_cnt_1_0_data_tmp[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_0));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[9].genblk1.PWM_int_RNO[9]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[9]), .C(
        un1_period_cnt_1_0), .Y(\un1_pwm_enable_reg_1_i_0[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[100]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[99]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[58]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[57]), .FCI(\un1_period_cnt_1_0_data_tmp_6[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_6[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[78]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[77]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[6] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f0[8]  (.A(
        \PWM_int_108_f1_14[8] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[8]), .D(\PWM_int_108_f1_13[8] ), .Y(
        \PWM_int_108[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[72]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[71]), .FCI(\un1_period_cnt_1_0_data_tmp_3[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_10[8]  (.A(
        pwm_negedge_reg[128]), .B(pwm_negedge_reg[122]), .C(
        pwm_negedge_reg[121]), .D(pwm_negedge_reg[120]), .Y(
        \PWM_int_108_f1_10[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[70]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[69]), .FCI(\un1_period_cnt_1_0_data_tmp_3[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[2] ));
    CFG4 #( .INIT(16'hC080) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0[3]  (.A(
        \PWM_int_38_f1_14[3] ), .B(un1_period_cnt_NE_i_0), .C(
        pwm_enable_reg[3]), .D(\PWM_int_38_f1_13[3] ), .Y(
        \PWM_int_38[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[126]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[125]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[6]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[5]), .FCI(\un1_period_cnt_1_0_data_tmp_1[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[26]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[25]), .FCI(\un1_period_cnt_1_0_data_tmp_0[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_0[4] ));
    SLE \PWM_output_generation[4].genblk1.PWM_int[4]  (.D(
        \PWM_int_52[4] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_8_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[4]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[138]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[137]), .FCI(
        \un1_period_cnt_1_0_data_tmp[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[4] ));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[4].genblk1.PWM_int_RNO[4]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[4]), .C(
        un1_period_cnt_1_7), .Y(\un1_pwm_enable_reg_8_i_0[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_3_4[5]  (.A(
        period_cnt[11]), .B(period_cnt[10]), .C(period_cnt[9]), .D(
        period_cnt[8]), .Y(\PWM_int_66_f0_i_3_4[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[80]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[79]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_4));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[56]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[55]), .FCI(\un1_period_cnt_1_0_data_tmp_6[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_6[3] ));
    CFG4 #( .INIT(16'h1333) )  
        \PWM_output_generation[7].genblk1.PWM_int_RNO[7]  (.A(
        \PWM_int_94_f0_i_a9_14[7] ), .B(\PWM_int_94_f0_i_1[7] ), .C(
        \PWM_int_94_f0_i_a9_10[7] ), .D(\PWM_int_94_f0_i_a9_9[7] ), .Y(
        N_29_i_0));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_39  (
        .A(pwm_negedge_reg[148]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[147]), .FCI(
        \un1_period_cnt_1_1_data_tmp[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[94]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[93]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[64]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[63]), .FCI(
        \un1_period_cnt_1_0_data_tmp_6[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_7));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f1_13[1]  (.A(
        pwm_negedge_reg[15]), .B(pwm_negedge_reg[16]), .C(
        \PWM_int_10_f1_10[1] ), .D(\PWM_int_10_f1_2[1] ), .Y(
        \PWM_int_10_f1_13[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[2]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[1]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[24]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[23]), .FCI(\un1_period_cnt_1_0_data_tmp_0[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_0[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[10].genblk1.un1_period_cnt_1_1_I_21  (
        .A(pwm_negedge_reg[152]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[151]), .FCI(
        \un1_period_cnt_1_1_data_tmp[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[136]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[135]), .FCI(
        \un1_period_cnt_1_0_data_tmp[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_3[5]  (.A(
        period_cnt[14]), .B(period_cnt[15]), .C(
        \PWM_int_66_f0_i_3_4[5] ), .D(\PWM_int_66_f0_i_3_3[5] ), .Y(
        N_29_3));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_8[3]  (.A(
        pwm_negedge_reg[42]), .B(pwm_negedge_reg[33]), .C(PWM_c[3]), 
        .Y(\PWM_int_38_f1_8[3] ));
    SLE \PWM_output_generation[8].genblk1.PWM_int[8]  (.D(
        \PWM_int_108[8] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_4_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[8]));
    CFG3 #( .INIT(8'hFB) )  
        \PWM_output_generation[6].genblk1.PWM_int_RNO[6]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[6]), .C(
        un1_period_cnt_1_3), .Y(\un1_pwm_enable_reg_2_i_0[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f1_10[3]  (.A(
        pwm_negedge_reg[48]), .B(pwm_negedge_reg[46]), .C(
        pwm_negedge_reg[45]), .D(pwm_negedge_reg[44]), .Y(
        \PWM_int_38_f1_10[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[122]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[121]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[4] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f1_2[2]  (.A(
        pwm_negedge_reg[27]), .B(pwm_negedge_reg[28]), .Y(
        \PWM_int_24_f1_2[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[12]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[11]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[5] ));
    CFG3 #( .INIT(8'hFB) )  \un1_pwm_enable_reg_3_i_0[0]  (.A(
        un1_period_cnt_NE_i_0), .B(pwm_enable_reg[5]), .C(
        un1_period_cnt_1_4), .Y(N_7));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[9].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[130]), .B(period_cnt[0]), .C(period_cnt[1]), 
        .D(pwm_negedge_reg[129]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[0] ));
    
endmodule


module timebase_16s(
       period_cnt,
       period_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST
    );
output [15:0] period_cnt;
input  [15:0] period_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;

    wire VCC_net_1, \period_cnt_s[0] , GND_net_1, \period_cnt_s[1] , 
        \period_cnt_s[2] , \period_cnt_s[3] , \period_cnt_s[4] , 
        \period_cnt_s[5] , \period_cnt_s[6] , \period_cnt_s[7] , 
        \period_cnt_s[8] , \period_cnt_s[9] , \period_cnt_s[10] , 
        \period_cnt_s[11] , \period_cnt_s[12] , \period_cnt_s[13] , 
        \period_cnt_s[14] , \period_cnt_s[15]_net_1 , 
        un1_period_cnt_cry_0_net_1, un1_period_cnt_cry_1_net_1, 
        un1_period_cnt_cry_2_net_1, un1_period_cnt_cry_3_net_1, 
        un1_period_cnt_cry_4_net_1, un1_period_cnt_cry_5_net_1, 
        un1_period_cnt_cry_6_net_1, un1_period_cnt_cry_7_net_1, 
        un1_period_cnt_cry_8_net_1, un1_period_cnt_cry_9_net_1, 
        un1_period_cnt_cry_10_net_1, un1_period_cnt_cry_11_net_1, 
        un1_period_cnt_cry_12_net_1, un1_period_cnt_cry_13_net_1, 
        un1_period_cnt_cry_14_net_1, period_cnt_net_1, 
        period_cnt_s_133_FCO, \period_cnt_cry[0]_net_1 , 
        \period_cnt_cry[1]_net_1 , \period_cnt_cry[2]_net_1 , 
        \period_cnt_cry[3]_net_1 , \period_cnt_cry[4]_net_1 , 
        \period_cnt_cry[5]_net_1 , \period_cnt_cry[6]_net_1 , 
        \period_cnt_cry[7]_net_1 , \period_cnt_cry[8]_net_1 , 
        \period_cnt_cry[9]_net_1 , \period_cnt_cry[10]_net_1 , 
        \period_cnt_cry[11]_net_1 , \period_cnt_cry[12]_net_1 , 
        \period_cnt_cry[13]_net_1 , \period_cnt_cry[14]_net_1 ;
    
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_9 (.A(period_reg[9])
        , .B(period_cnt[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_8_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_9_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_2 (.A(period_reg[2])
        , .B(period_cnt[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_1_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_2_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[14]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[14]), .D(GND_net_1), .FCI(
        \period_cnt_cry[13]_net_1 ), .S(\period_cnt_s[14] ), .Y(), 
        .FCO(\period_cnt_cry[14]_net_1 ));
    SLE \period_cnt[9]  (.D(\period_cnt_s[9] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[9]));
    SLE \period_cnt[6]  (.D(\period_cnt_s[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[6]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[0]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[0]), .D(GND_net_1), .FCI(
        period_cnt_s_133_FCO), .S(\period_cnt_s[0] ), .Y(), .FCO(
        \period_cnt_cry[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  period_cnt_s_133 (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(period_cnt_s_133_FCO));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[8]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[8]), .D(GND_net_1), .FCI(
        \period_cnt_cry[7]_net_1 ), .S(\period_cnt_s[8] ), .Y(), .FCO(
        \period_cnt_cry[8]_net_1 ));
    SLE \period_cnt[14]  (.D(\period_cnt_s[14] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[14]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[11]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[11]), .D(GND_net_1), .FCI(
        \period_cnt_cry[10]_net_1 ), .S(\period_cnt_s[11] ), .Y(), 
        .FCO(\period_cnt_cry[11]_net_1 ));
    SLE \period_cnt[10]  (.D(\period_cnt_s[10] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[10]));
    SLE \period_cnt[0]  (.D(\period_cnt_s[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[0]));
    SLE \period_cnt[11]  (.D(\period_cnt_s[11] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[11]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_3 (.A(period_reg[3])
        , .B(period_cnt[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_2_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_3_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE \period_cnt[13]  (.D(\period_cnt_s[13] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[13]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[7]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[7]), .D(GND_net_1), .FCI(
        \period_cnt_cry[6]_net_1 ), .S(\period_cnt_s[7] ), .Y(), .FCO(
        \period_cnt_cry[7]_net_1 ));
    SLE \period_cnt[1]  (.D(\period_cnt_s[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[1]));
    SLE \period_cnt[7]  (.D(\period_cnt_s[7] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[7]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[1]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[1]), .D(GND_net_1), .FCI(
        \period_cnt_cry[0]_net_1 ), .S(\period_cnt_s[1] ), .Y(), .FCO(
        \period_cnt_cry[1]_net_1 ));
    SLE \period_cnt[15]  (.D(\period_cnt_s[15]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(period_cnt[15]));
    SLE \period_cnt[2]  (.D(\period_cnt_s[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[2]));
    SLE \period_cnt[3]  (.D(\period_cnt_s[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[3]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_5 (.A(period_reg[5])
        , .B(period_cnt[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_4_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_5_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[9]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[9]), .D(GND_net_1), .FCI(
        \period_cnt_cry[8]_net_1 ), .S(\period_cnt_s[9] ), .Y(), .FCO(
        \period_cnt_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[2]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[2]), .D(GND_net_1), .FCI(
        \period_cnt_cry[1]_net_1 ), .S(\period_cnt_s[2] ), .Y(), .FCO(
        \period_cnt_cry[2]_net_1 ));
    SLE \period_cnt[5]  (.D(\period_cnt_s[5] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[5]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_11 (.A(
        period_reg[11]), .B(period_cnt[11]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_10_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_11_net_1));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[10]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[10]), .D(GND_net_1), .FCI(
        \period_cnt_cry[9]_net_1 ), .S(\period_cnt_s[10] ), .Y(), .FCO(
        \period_cnt_cry[10]_net_1 ));
    SLE \period_cnt[4]  (.D(\period_cnt_s[4] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[4]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_8 (.A(period_reg[8])
        , .B(period_cnt[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_7_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_8_net_1));
    SLE \period_cnt[8]  (.D(\period_cnt_s[8] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[8]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_10 (.A(
        period_reg[10]), .B(period_cnt[10]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_9_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_10_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[12]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[12]), .D(GND_net_1), .FCI(
        \period_cnt_cry[11]_net_1 ), .S(\period_cnt_s[12] ), .Y(), 
        .FCO(\period_cnt_cry[12]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_4 (.A(period_reg[4])
        , .B(period_cnt[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_3_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_4_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_14 (.A(
        period_reg[14]), .B(period_cnt[14]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_13_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_14_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_7 (.A(period_reg[7])
        , .B(period_cnt[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_6_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_7_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_15 (.A(
        period_reg[15]), .B(period_cnt[15]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_14_net_1), .S(), .Y(), 
        .FCO(period_cnt_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[3]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[3]), .D(GND_net_1), .FCI(
        \period_cnt_cry[2]_net_1 ), .S(\period_cnt_s[3] ), .Y(), .FCO(
        \period_cnt_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[5]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[5]), .D(GND_net_1), .FCI(
        \period_cnt_cry[4]_net_1 ), .S(\period_cnt_s[5] ), .Y(), .FCO(
        \period_cnt_cry[5]_net_1 ));
    SLE \period_cnt[12]  (.D(\period_cnt_s[12] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[12]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_0 (.A(period_reg[0])
        , .B(period_cnt[0]), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(un1_period_cnt_cry_0_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[4]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[4]), .D(GND_net_1), .FCI(
        \period_cnt_cry[3]_net_1 ), .S(\period_cnt_s[4] ), .Y(), .FCO(
        \period_cnt_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_6 (.A(period_reg[6])
        , .B(period_cnt[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_5_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_6_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_12 (.A(
        period_reg[12]), .B(period_cnt[12]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_11_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_12_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_1 (.A(period_reg[1])
        , .B(period_cnt[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_0_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_1_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_s[15]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[15]), .D(GND_net_1), .FCI(
        \period_cnt_cry[14]_net_1 ), .S(\period_cnt_s[15]_net_1 ), .Y()
        , .FCO());
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_13 (.A(
        period_reg[13]), .B(period_cnt[13]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_12_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_13_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[13]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[13]), .D(GND_net_1), .FCI(
        \period_cnt_cry[12]_net_1 ), .S(\period_cnt_s[13] ), .Y(), 
        .FCO(\period_cnt_cry[13]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[6]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[6]), .D(GND_net_1), .FCI(
        \period_cnt_cry[5]_net_1 ), .S(\period_cnt_s[6] ), .Y(), .FCO(
        \period_cnt_cry[6]_net_1 ));
    
endmodule


module reg_if_Z6(
       CoreAPB3_0_APBmslave0_PWDATA,
       pwm_enable_reg,
       pwm_negedge_reg,
       period_reg,
       period_cnt,
       iPSELS_0_0,
       iPSELS_0,
       CoreAPB3_0_APBmslave0_PADDR,
       CoreAPB3_0_APBmslave4_PRDATA,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       N_97_1,
       controlReg14_3,
       PRDATA_regif_sn_N_26,
       N_842,
       N_841,
       N_840,
       un1_OEn_2,
       un3_PRDATA_regif_1,
       psh_negedge_reg_1_sqmuxa_3_2,
       N_813,
       N_811,
       N_806,
       N_812,
       N_807,
       N_808,
       N_810,
       N_809,
       controlReg24_3,
       PRDATA_regif_sn_N_39_mux,
       N_833,
       N_831,
       N_828,
       N_826,
       N_832,
       N_827,
       N_830,
       N_829,
       N_837,
       N_839,
       N_838
    );
input  [15:0] CoreAPB3_0_APBmslave0_PWDATA;
output [10:1] pwm_enable_reg;
output [160:1] pwm_negedge_reg;
output [15:0] period_reg;
input  [15:0] period_cnt;
input  [4:4] iPSELS_0_0;
input  [4:4] iPSELS_0;
input  [7:2] CoreAPB3_0_APBmslave0_PADDR;
output [1:0] CoreAPB3_0_APBmslave4_PRDATA;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  N_97_1;
input  controlReg14_3;
output PRDATA_regif_sn_N_26;
output N_842;
output N_841;
output N_840;
input  un1_OEn_2;
output un3_PRDATA_regif_1;
output psh_negedge_reg_1_sqmuxa_3_2;
output N_813;
output N_811;
output N_806;
output N_812;
output N_807;
output N_808;
output N_810;
output N_809;
input  controlReg24_3;
output PRDATA_regif_sn_N_39_mux;
output N_833;
output N_831;
output N_828;
output N_826;
output N_832;
output N_827;
output N_830;
output N_829;
output N_837;
output N_839;
output N_838;

    wire un1_period_cnt, un1_period_cnt_i_0, VCC_net_1, 
        psh_negedge_reg_1_sqmuxa_1_net_1, GND_net_1, 
        psh_negedge_reg_1_sqmuxa_net_1, 
        psh_negedge_reg_1_sqmuxa_7_net_1, 
        psh_negedge_reg_1_sqmuxa_3_net_1, 
        psh_enable_reg1_1_sqmuxa_net_1, psh_enable_reg2_1_sqmuxa_net_1, 
        psh_negedge_reg_1_sqmuxa_6_net_1, 
        psh_negedge_reg_1_sqmuxa_9_net_1, 
        psh_negedge_reg_1_sqmuxa_5_net_1, 
        psh_negedge_reg_1_sqmuxa_4_net_1, 
        psh_negedge_reg_1_sqmuxa_8_net_1, 
        psh_negedge_reg_1_sqmuxa_2_net_1, \psh_period_reg[4]_net_1 , 
        \psh_period_reg[5]_net_1 , \psh_period_reg[6]_net_1 , 
        \psh_period_reg[7]_net_1 , \psh_period_reg[8]_net_1 , 
        \psh_period_reg[9]_net_1 , \psh_period_reg[10]_net_1 , 
        \psh_period_reg[11]_net_1 , \psh_period_reg[12]_net_1 , 
        \psh_period_reg[13]_net_1 , \psh_period_reg[14]_net_1 , 
        \psh_period_reg[15]_net_1 , psh_period_reg_1_sqmuxa_net_1, 
        \psh_period_reg[0]_net_1 , \psh_period_reg[1]_net_1 , 
        \psh_period_reg[2]_net_1 , \psh_period_reg[3]_net_1 , 
        sync_update_net_1, sync_update_0_sqmuxa_net_1, 
        un1_period_cnt_cry_0, un1_period_cnt_cry_1, 
        un1_period_cnt_cry_2, un1_period_cnt_cry_3, 
        un1_period_cnt_cry_4, un1_period_cnt_cry_5, 
        un1_period_cnt_cry_6, un1_period_cnt_cry_7, 
        un1_period_cnt_cry_8, un1_period_cnt_cry_9, 
        un1_period_cnt_cry_10, un1_period_cnt_cry_11, 
        un1_period_cnt_cry_12, un1_period_cnt_cry_13, 
        un1_period_cnt_cry_14, psh_prescale_reg13_net_1, 
        PRDATA_regif_13_N_2L1_net_1, PRDATA_regif_sn_m21_a1_1_net_1, 
        PRDATA_regif_13_N_4L5_net_1, PRDATA_regif_sn_m21_a0_0_net_1, 
        PRDATA_regif_13_N_5L8_net_1, N_762, N_815, 
        \PRDATA_regif_15_am_1[7]_net_1 , 
        \PRDATA_regif_15_am_1_0[7]_net_1 , 
        \PRDATA_regif_15_am[7]_net_1 , \PRDATA_regif_15_am_1[6]_net_1 , 
        \PRDATA_regif_15_am_1_0[6]_net_1 , 
        \PRDATA_regif_15_am[6]_net_1 , \PRDATA_regif_15_am_1[5]_net_1 , 
        \PRDATA_regif_15_am_1_0[5]_net_1 , 
        \PRDATA_regif_15_am[5]_net_1 , PRDATA_regif_sn_m25_1_net_1, 
        \PRDATA_regif_12_1[1] , \PRDATA_regif_12_1_0[1] , N_799, 
        \PRDATA_regif_12_1[4] , \PRDATA_regif_12_1_0[4] , N_802, 
        \PRDATA_regif_12_1[2] , \PRDATA_regif_12_1_0[2] , N_800, 
        \PRDATA_regif_12_1[0] , \PRDATA_regif_12_1_0[0] , N_798, 
        \PRDATA_regif_12_1[3] , \PRDATA_regif_12_1_0[3] , N_801, 
        \PRDATA_regif_10_1_1[9] , N_773, \PRDATA_regif_10_1_1[4] , 
        N_768, \PRDATA_regif_10_1[0] , N_764, 
        \PRDATA_regif_10_1_1[14] , N_778, \PRDATA_regif_10_1_1[11] , 
        N_775, \PRDATA_regif_10_1_1[3] , N_767, 
        \PRDATA_regif_10_1_1[8] , N_772, \PRDATA_regif_10_1_1[12] , 
        N_776, \PRDATA_regif_10_1_1[10] , N_774, 
        \PRDATA_regif_10_1[1] , N_765, \PRDATA_regif_10_1_1[6] , N_770, 
        \PRDATA_regif_10_1_1[7] , N_771, \PRDATA_regif_10_1_1[13] , 
        N_777, \PRDATA_regif_10_1_1[15] , N_779, 
        \PRDATA_regif_10_1_1[5] , N_769, \PRDATA_regif_10_1_1[2] , 
        N_766, \PRDATA_regif_15_bm[7]_net_1 , 
        \PRDATA_regif_15_bm[6]_net_1 , \PRDATA_regif_15_bm[5]_net_1 , 
        \PRDATA_regif_11_bm[1]_net_1 , \PRDATA_regif_11_am[1]_net_1 , 
        N_781, \PRDATA_regif_11_bm[11]_net_1 , 
        \PRDATA_regif_11_am[11]_net_1 , N_791, 
        \PRDATA_regif_11_bm[12]_net_1 , \PRDATA_regif_11_am[12]_net_1 , 
        N_792, \PRDATA_regif_11_bm[9]_net_1 , 
        \PRDATA_regif_11_am[9]_net_1 , N_789, 
        \PRDATA_regif_11_bm[7]_net_1 , \PRDATA_regif_11_am[7]_net_1 , 
        N_787, \PRDATA_regif_11_bm[14]_net_1 , 
        \PRDATA_regif_11_am[14]_net_1 , N_794, 
        \PRDATA_regif_11_bm[0]_net_1 , \PRDATA_regif_11_am[0]_net_1 , 
        N_780, \PRDATA_regif_11_bm[3]_net_1 , 
        \PRDATA_regif_11_am[3]_net_1 , N_783, 
        \PRDATA_regif_11_bm[2]_net_1 , \PRDATA_regif_11_am[2]_net_1 , 
        N_782, \PRDATA_regif_11_bm[5]_net_1 , 
        \PRDATA_regif_11_am[5]_net_1 , N_785, 
        \PRDATA_regif_11_bm[6]_net_1 , \PRDATA_regif_11_am[6]_net_1 , 
        N_786, \PRDATA_regif_11_bm[8]_net_1 , 
        \PRDATA_regif_11_am[8]_net_1 , N_788, 
        \PRDATA_regif_11_bm[4]_net_1 , \PRDATA_regif_11_am[4]_net_1 , 
        N_784, \PRDATA_regif_11_bm[10]_net_1 , 
        \PRDATA_regif_11_am[10]_net_1 , N_790, 
        \PRDATA_regif_11_bm[13]_net_1 , \PRDATA_regif_11_am[13]_net_1 , 
        N_793, \PRDATA_regif_11_bm[15]_net_1 , 
        \PRDATA_regif_11_am[15]_net_1 , N_795, 
        \PRDATA_regif_13_1[1]_net_1 , N_816, 
        psh_negedge_reg_1_sqmuxa_8_1_net_1, 
        psh_negedge_reg_1_sqmuxa_5_2, N_743, N_741, N_736, N_742, 
        PRDATA_regif_sn_N_15, N_737, N_738, N_740, N_739, 
        psh_enable_reg1_1_sqmuxa_2_net_1, 
        psh_negedge_reg_1_sqmuxa_4_1_net_1, 
        psh_negedge_reg_1_sqmuxa_1_1_net_1, 
        psh_negedge_reg_1_sqmuxa_1_0_net_1, 
        psh_period_reg_1_sqmuxa_1_net_1, 
        psh_negedge_reg_1_sqmuxa_6_1_net_1, 
        psh_negedge_reg_1_sqmuxa_7_1_net_1, 
        psh_negedge_reg_1_sqmuxa_8_1_0, sync_update_0_sqmuxa_1_net_1, 
        psh_negedge_reg_1_sqmuxa_3_0_net_1, 
        \PRDATA_regif_9_1[0]_net_1 , 
        psh_enable_reg2_1_sqmuxa_1_0_net_1, N_822, N_820, N_821, N_818, 
        N_819, N_835, N_836;
    
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[14]  (.A(
        pwm_negedge_reg[143]), .B(pwm_negedge_reg[95]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_742));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[70]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[70]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[42]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[42]));
    CFG2 #( .INIT(4'h7) )  PRDATA_regif_13_N_4L5 (.A(
        PRDATA_regif_sn_m21_a1_1_net_1), .B(N_97_1), .Y(
        PRDATA_regif_13_N_4L5_net_1));
    SLE \period_reg[5]  (.D(\psh_period_reg[5]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[5]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[27]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[27]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[126]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[126]));
    SLE \period_reg[14]  (.D(\psh_period_reg[14]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[14]));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[13]  (.A(
        pwm_negedge_reg[46]), .B(pwm_negedge_reg[110]), .C(
        \PRDATA_regif_10_1_1[13] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_777));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[111]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[111]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_1[3]  (.A(
        pwm_negedge_reg[84]), .B(pwm_enable_reg[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\PRDATA_regif_12_1_0[3] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_15  (.A(period_reg[15])
        , .B(period_cnt[15]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_14), .S(), .Y(), .FCO(un1_period_cnt));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[14]  (.A(
        pwm_negedge_reg[47]), .B(pwm_negedge_reg[111]), .C(
        \PRDATA_regif_10_1_1[14] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_778));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[45]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[45]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[150]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[150]));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[8]  (.A(
        pwm_negedge_reg[137]), .B(pwm_negedge_reg[89]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_736));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[131]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[131]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[14]  (.A(
        pwm_negedge_reg[79]), .B(pwm_negedge_reg[15]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[14]_net_1 ));
    SLE \period_reg[12]  (.D(\psh_period_reg[12]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[12]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_8  (.A(period_reg[8]), 
        .B(period_cnt[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_7), .S(), .Y(), .FCO(un1_period_cnt_cry_8));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_15_bm_RNO[5]  (.A(
        pwm_negedge_reg[38]), .B(pwm_negedge_reg[102]), .C(
        \PRDATA_regif_10_1_1[5] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_769));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[82]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[82]));
    SLE \psh_period_reg[14]  (.D(CoreAPB3_0_APBmslave0_PWDATA[14]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[14]_net_1 )
        );
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_1[4]  (.A(
        pwm_negedge_reg[85]), .B(pwm_enable_reg[5]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\PRDATA_regif_12_1_0[4] ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[89]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[89]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[57]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[57]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[69]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[69]));
    CFG4 #( .INIT(16'h2000) )  psh_negedge_reg_1_sqmuxa_3 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        psh_negedge_reg_1_sqmuxa_3_0_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_3_net_1)
        );
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[79]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[79]));
    SLE \period_reg[13]  (.D(\psh_period_reg[13]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[13]));
    CFG4 #( .INIT(16'h1000) )  psh_negedge_reg_1_sqmuxa_4 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_negedge_reg_1_sqmuxa_4_1_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_4_net_1)
        );
    SLE \period_reg[8]  (.D(\psh_period_reg[8]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[8]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[101]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[101]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[20]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[20]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[153]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[153]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[157]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[157]));
    CFG3 #( .INIT(8'h1B) )  PRDATA_regif_sn_m14 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(PRDATA_regif_sn_N_15));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_15_bm_RNO_0[7]  (.A(
        pwm_negedge_reg[56]), .B(pwm_negedge_reg[120]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[7] ));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[135]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[135]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_1[1]  (.A(
        pwm_negedge_reg[82]), .B(pwm_enable_reg[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\PRDATA_regif_12_1_0[1] ));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[141]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[141]));
    SLE \period_reg[11]  (.D(\psh_period_reg[11]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[11]));
    SLE \psh_period_reg[12]  (.D(CoreAPB3_0_APBmslave0_PWDATA[12]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[12]_net_1 )
        );
    SLE \psh_enable_reg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[4]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[92]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[92]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[97]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[97]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1_0[6]  (.A(
        pwm_negedge_reg[87]), .B(pwm_enable_reg[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_regif_15_am_1_0[6]_net_1 ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[37]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[37]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[136]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[136]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[8]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[8]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[23]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[23]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[1]  (.A(
        pwm_negedge_reg[50]), .B(pwm_negedge_reg[114]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1[1] ));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[11]  (.A(
        pwm_negedge_reg[44]), .B(pwm_negedge_reg[108]), .C(
        \PRDATA_regif_10_1_1[11] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_775));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[9]  (.A(
        pwm_negedge_reg[74]), .B(pwm_negedge_reg[10]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[9]_net_1 ));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[149]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[149]));
    SLE \period_reg[3]  (.D(\psh_period_reg[3]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[3]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[65]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[65]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[119]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[119]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[105]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[105]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[154]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[154]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[1]  (.A(
        pwm_negedge_reg[146]), .B(pwm_negedge_reg[18]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[1]_net_1 ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[46]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[46]));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[4]  (.A(
        pwm_negedge_reg[37]), .B(pwm_negedge_reg[101]), .C(
        \PRDATA_regif_10_1_1[4] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_768));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[75]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[75]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[2]  (.A(
        pwm_negedge_reg[147]), .B(pwm_negedge_reg[19]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[2]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[9]  (.A(N_773), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_789), .Y(N_827));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_14  (.A(period_reg[14])
        , .B(period_cnt[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_13), .S(), .Y(), .FCO(un1_period_cnt_cry_14)
        );
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[106]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[106]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[35]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[35]));
    SLE \psh_period_reg[8]  (.D(CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[8]_net_1 ));
    SLE \period_reg[0]  (.D(\psh_period_reg[0]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[0]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_15_bm[6]  (.A(N_770), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_786), .Y(
        \PRDATA_regif_15_bm[6]_net_1 ));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_15_bm_RNO[7]  (.A(
        pwm_negedge_reg[40]), .B(pwm_negedge_reg[104]), .C(
        \PRDATA_regif_10_1_1[7] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_771));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[0]  (.A(
        \PRDATA_regif_11_bm[0]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[0]_net_1 ), .Y(N_780));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[14]  (.A(N_742), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[14]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_812));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[58]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[58]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[12]  (.A(N_776), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_792), .Y(N_830));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[2]  (.A(N_766), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_782), .Y(N_820));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[10]  (.A(N_738), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[10]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_808));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[7]  (.A(
        pwm_negedge_reg[152]), .B(pwm_negedge_reg[24]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[7]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[114]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[114]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[60]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[60]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[44]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[44]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_0[4]  (.A(
        pwm_negedge_reg[133]), .B(period_reg[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\PRDATA_regif_12_1[4] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_1  (.A(period_reg[1]), 
        .B(period_cnt[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_0), .S(), .Y(), .FCO(un1_period_cnt_cry_1));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[0]  (.A(
        pwm_negedge_reg[65]), .B(pwm_negedge_reg[1]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[0]_net_1 ));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_am[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        \PRDATA_regif_15_am_1[7]_net_1 ), .C(
        \PRDATA_regif_15_am_1_0[7]_net_1 ), .Y(
        \PRDATA_regif_15_am[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_15_RNIHOI2  (.A(
        un1_period_cnt), .Y(un1_period_cnt_i_0));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[4]  (.A(
        \PRDATA_regif_11_bm[4]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[4]_net_1 ), .Y(N_784));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[118]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[118]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[87]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[87]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_11  (.A(period_reg[11])
        , .B(period_cnt[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_10), .S(), .Y(), .FCO(un1_period_cnt_cry_11)
        );
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[5]  (.A(
        pwm_negedge_reg[70]), .B(pwm_negedge_reg[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[5]_net_1 ));
    SLE \psh_period_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[2]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[80]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[80]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[147]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[147]));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[13]  (.A(N_741), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[13]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_811));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[68]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[68]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[62]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[62]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[10]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[10]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[12]  (.A(
        pwm_negedge_reg[157]), .B(pwm_negedge_reg[29]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[12]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[78]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[78]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[15]  (.A(
        pwm_negedge_reg[80]), .B(pwm_negedge_reg[16]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[15]_net_1 ));
    SLE \psh_period_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[1]_net_1 ));
    CFG2 #( .INIT(4'h2) )  psh_negedge_reg_1_sqmuxa_2_3 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        psh_negedge_reg_1_sqmuxa_5_2));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1[7]  (.A(
        pwm_negedge_reg[136]), .B(period_reg[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_15_am_1[7]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[1]  (.A(N_765), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_781), .Y(N_819));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15_ns[5]  (.A(
        \PRDATA_regif_15_bm[5]_net_1 ), .B(
        \PRDATA_regif_15_am[5]_net_1 ), .C(PRDATA_regif_sn_N_26), .Y(
        N_840));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[12]  (.A(
        pwm_negedge_reg[61]), .B(pwm_negedge_reg[125]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[12] ));
    SLE \psh_period_reg[10]  (.D(CoreAPB3_0_APBmslave0_PWDATA[10]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[10]_net_1 )
        );
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[8]  (.A(
        pwm_negedge_reg[153]), .B(pwm_negedge_reg[25]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[8]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[3]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[3]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[13]  (.A(
        pwm_negedge_reg[78]), .B(pwm_negedge_reg[14]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[13]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[4]  (.A(
        pwm_negedge_reg[69]), .B(pwm_negedge_reg[5]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[4]_net_1 ));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[127]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[127]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[28]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[28]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[36]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[36]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_7  (.A(period_reg[7]), 
        .B(period_cnt[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_6), .S(), .Y(), .FCO(un1_period_cnt_cry_7));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_0[3]  (.A(
        pwm_negedge_reg[132]), .B(period_reg[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\PRDATA_regif_12_1[3] ));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[22]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[22]));
    CFG4 #( .INIT(16'h0008) )  psh_negedge_reg_1_sqmuxa_6_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        psh_negedge_reg_1_sqmuxa_6_1_net_1));
    CFG3 #( .INIT(8'h20) )  sync_update_0_sqmuxa (.A(
        psh_prescale_reg13_net_1), .B(un3_PRDATA_regif_1), .C(
        sync_update_0_sqmuxa_1_net_1), .Y(sync_update_0_sqmuxa_net_1));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[11]  (.A(
        \PRDATA_regif_11_bm[11]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[11]_net_1 ), .Y(N_791));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_RNO[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\PRDATA_regif_12_1[4] ), 
        .C(\PRDATA_regif_12_1_0[4] ), .Y(N_802));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[8]  (.A(
        pwm_negedge_reg[57]), .B(pwm_negedge_reg[121]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[8] ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[11]  (.A(
        pwm_negedge_reg[76]), .B(pwm_negedge_reg[12]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[11]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[15]  (.A(
        \PRDATA_regif_11_bm[15]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[15]_net_1 ), .Y(N_795));
    SLE \psh_period_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[15]  (.A(N_779), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_795), .Y(N_833));
    CFG2 #( .INIT(4'h7) )  PRDATA_regif_13_N_2L1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(sync_update_net_1), .Y(
        PRDATA_regif_13_N_2L1_net_1));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[15]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[15]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[84]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[84]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[3]  (.A(
        pwm_negedge_reg[52]), .B(pwm_negedge_reg[116]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[3] ));
    CFG4 #( .INIT(16'h8B0F) )  \PRDATA_regif_13[0]  (.A(N_762), .B(
        PRDATA_regif_13_N_5L8_net_1), .C(PRDATA_regif_13_N_2L1_net_1), 
        .D(PRDATA_regif_13_N_4L5_net_1), .Y(N_815));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[4]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[4]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[34]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[34]));
    CFG4 #( .INIT(16'h7000) )  \PRDATA_regif_13_1[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(pwm_enable_reg[10]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_regif_13_1[1]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \PRDATA_regif_13[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[7]), .B(un1_OEn_2), .C(
        \PRDATA_regif_13_1[1]_net_1 ), .Y(N_816));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[10]  (.A(
        pwm_negedge_reg[43]), .B(pwm_negedge_reg[107]), .C(
        \PRDATA_regif_10_1_1[10] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_774));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15_ns[7]  (.A(
        \PRDATA_regif_15_bm[7]_net_1 ), .B(
        \PRDATA_regif_15_am[7]_net_1 ), .C(PRDATA_regif_sn_N_26), .Y(
        N_842));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[13]  (.A(
        \PRDATA_regif_11_bm[13]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[13]_net_1 ), .Y(N_793));
    SLE \period_reg[9]  (.D(\psh_period_reg[9]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[9]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[123]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[123]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[5]  (.A(
        \PRDATA_regif_11_bm[5]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[5]_net_1 ), .Y(N_785));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[50]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[50]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[14]  (.A(
        \PRDATA_regif_11_bm[14]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[14]_net_1 ), .Y(N_794));
    SLE \period_reg[2]  (.D(\psh_period_reg[2]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[2]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15[3]  (.A(N_821), .B(N_801), 
        .C(PRDATA_regif_sn_N_26), .Y(N_838));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_3  (.A(period_reg[3]), 
        .B(period_cnt[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_2), .S(), .Y(), .FCO(un1_period_cnt_cry_3));
    CFG4 #( .INIT(16'h8000) )  sync_update_0_sqmuxa_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        sync_update_0_sqmuxa_1_net_1));
    SLE \psh_period_reg[13]  (.D(CoreAPB3_0_APBmslave0_PWDATA[13]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[13]_net_1 )
        );
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[10]  (.A(
        pwm_negedge_reg[155]), .B(pwm_negedge_reg[27]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[10]_net_1 ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[94]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[94]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[137]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[137]));
    SLE \psh_enable_reg1[8]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[8]));
    CFG4 #( .INIT(16'hB8AA) )  \PRDATA_regif[1]  (.A(N_816), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(N_836), .D(
        PRDATA_regif_sn_N_39_mux), .Y(CoreAPB3_0_APBmslave4_PRDATA[1]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[151]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[151]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_15_bm_RNO_0[6]  (.A(
        pwm_negedge_reg[55]), .B(pwm_negedge_reg[119]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[6] ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15[2]  (.A(N_820), .B(N_800), 
        .C(PRDATA_regif_sn_N_26), .Y(N_837));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[52]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[52]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[31]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[31]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1_0[5]  (.A(
        pwm_negedge_reg[86]), .B(pwm_enable_reg[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_regif_15_am_1_0[5]_net_1 ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[40]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[40]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[1]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[1]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[12]  (.A(
        \PRDATA_regif_11_bm[12]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[12]_net_1 ), .Y(N_792));
    SLE \psh_period_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[5]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[0]  (.A(N_764), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_780), .Y(N_818));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[6]  (.A(
        pwm_negedge_reg[151]), .B(pwm_negedge_reg[23]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[6]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_4  (.A(period_reg[4]), 
        .B(period_cnt[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_3), .S(), .Y(), .FCO(un1_period_cnt_cry_4));
    SLE sync_update (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(sync_update_0_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(sync_update_net_1));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[1]  (.A(
        pwm_negedge_reg[66]), .B(pwm_negedge_reg[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[1]_net_1 ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[107]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[107]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[71]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[71]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[3]  (.A(
        pwm_negedge_reg[148]), .B(pwm_negedge_reg[20]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[12]  (.A(
        pwm_negedge_reg[77]), .B(pwm_negedge_reg[13]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[12]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[7]  (.A(
        \PRDATA_regif_11_bm[7]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[7]_net_1 ), .Y(N_787));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_am[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        \PRDATA_regif_15_am_1[6]_net_1 ), .C(
        \PRDATA_regif_15_am_1_0[6]_net_1 ), .Y(
        \PRDATA_regif_15_am[6]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[2]  (.A(
        pwm_negedge_reg[67]), .B(pwm_negedge_reg[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[2]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[10]  (.A(
        pwm_negedge_reg[75]), .B(pwm_negedge_reg[11]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[10]_net_1 ));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[115]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[115]));
    CFG4 #( .INIT(16'h0080) )  psh_negedge_reg_1_sqmuxa_7_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        psh_negedge_reg_1_sqmuxa_7_1_net_1));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15_ns[6]  (.A(
        \PRDATA_regif_15_bm[6]_net_1 ), .B(
        \PRDATA_regif_15_am[6]_net_1 ), .C(PRDATA_regif_sn_N_26), .Y(
        N_841));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[2]  (.A(
        pwm_negedge_reg[35]), .B(pwm_negedge_reg[99]), .C(
        \PRDATA_regif_10_1_1[2] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_766));
    SLE \period_reg[4]  (.D(\psh_period_reg[4]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[4]));
    CFG4 #( .INIT(16'h2000) )  psh_negedge_reg_1_sqmuxa_9 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_enable_reg2_1_sqmuxa_1_0_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_9_net_1)
        );
    CFG4 #( .INIT(16'hACAA) )  \PRDATA_regif[0]  (.A(N_815), .B(N_835), 
        .C(CoreAPB3_0_APBmslave0_PADDR[7]), .D(
        PRDATA_regif_sn_N_39_mux), .Y(CoreAPB3_0_APBmslave4_PRDATA[0]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[133]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[133]));
    CFG4 #( .INIT(16'h1000) )  psh_negedge_reg_1_sqmuxa (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_negedge_reg_1_sqmuxa_1_1_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_net_1));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[116]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[116]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[43]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[43]));
    CFG4 #( .INIT(16'h1000) )  psh_enable_reg1_1_sqmuxa (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_enable_reg1_1_sqmuxa_2_net_1), .D(psh_prescale_reg13_net_1)
        , .Y(psh_enable_reg1_1_sqmuxa_net_1));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15[0]  (.A(N_818), .B(N_798), 
        .C(PRDATA_regif_sn_N_26), .Y(N_835));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[7]  (.A(
        pwm_negedge_reg[72]), .B(pwm_negedge_reg[8]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[7]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \genblk1.un3_PRDATA_regiflto5_1  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(un3_PRDATA_regif_1));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[2]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[2]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1_0[7]  (.A(
        pwm_negedge_reg[88]), .B(pwm_enable_reg[8]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_regif_15_am_1_0[7]_net_1 ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[85]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[85]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_0[0]  (.A(
        pwm_negedge_reg[129]), .B(period_reg[0]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\PRDATA_regif_12_1[0] ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[9]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[9]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[14]  (.A(
        pwm_negedge_reg[159]), .B(pwm_negedge_reg[31]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[14]_net_1 ));
    CFG3 #( .INIT(8'h08) )  psh_negedge_reg_1_sqmuxa_3_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        psh_negedge_reg_1_sqmuxa_3_2), .C(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        psh_negedge_reg_1_sqmuxa_3_0_net_1));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[8]  (.A(N_772), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_788), .Y(N_826));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[1]  (.A(
        pwm_negedge_reg[34]), .B(pwm_negedge_reg[98]), .C(
        \PRDATA_regif_10_1[1] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_765));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[103]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[103]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[63]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[63]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[13]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[13]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15[4]  (.A(N_822), .B(N_802), 
        .C(PRDATA_regif_sn_N_26), .Y(N_839));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[12]  (.A(N_740), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[12]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_810));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[88]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[88]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1[6]  (.A(
        pwm_negedge_reg[135]), .B(period_reg[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_15_am_1[6]_net_1 ));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[143]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[143]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[64]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[64]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[73]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[73]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[155]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[155]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[11]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[11]));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[12]  (.A(
        pwm_negedge_reg[45]), .B(pwm_negedge_reg[109]), .C(
        \PRDATA_regif_10_1_1[12] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_776));
    CFG2 #( .INIT(4'h1) )  PRDATA_regif_sn_m21_a0_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[7]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        PRDATA_regif_sn_m21_a0_0_net_1));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[9]  (.A(
        pwm_negedge_reg[138]), .B(pwm_negedge_reg[90]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_737));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[10]  (.A(
        pwm_negedge_reg[139]), .B(pwm_negedge_reg[91]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_738));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[0]  (.A(
        pwm_negedge_reg[33]), .B(pwm_negedge_reg[97]), .C(
        \PRDATA_regif_10_1[0] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_764));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[120]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[120]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[3]  (.A(N_767), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_783), .Y(N_821));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[99]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[99]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[2]  (.A(
        pwm_negedge_reg[51]), .B(pwm_negedge_reg[115]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[2] ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[6]  (.A(
        \PRDATA_regif_11_bm[6]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[6]_net_1 ), .Y(N_786));
    CFG4 #( .INIT(16'h0800) )  PRDATA_regif_sn_m21_a1_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        PRDATA_regif_sn_m21_a1_1_net_1));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[95]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[95]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_2  (.A(period_reg[2]), 
        .B(period_cnt[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_1), .S(), .Y(), .FCO(un1_period_cnt_cry_2));
    SLE \psh_period_reg[11]  (.D(CoreAPB3_0_APBmslave0_PWDATA[11]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[11]_net_1 )
        );
    CFG4 #( .INIT(16'h0800) )  psh_negedge_reg_1_sqmuxa_1_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        psh_negedge_reg_1_sqmuxa_1_1_net_1));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[8]  (.A(
        \PRDATA_regif_11_bm[8]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[8]_net_1 ), .Y(N_788));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[8]  (.A(
        pwm_negedge_reg[73]), .B(pwm_negedge_reg[9]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[8]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_15[1]  (.A(N_819), .B(N_799), 
        .C(PRDATA_regif_sn_N_26), .Y(N_836));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_5  (.A(period_reg[5]), 
        .B(period_cnt[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_4), .S(), .Y(), .FCO(un1_period_cnt_cry_5));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_15_bm_RNO[6]  (.A(
        pwm_negedge_reg[39]), .B(pwm_negedge_reg[103]), .C(
        \PRDATA_regif_10_1_1[6] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_770));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[25]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[25]));
    CFG3 #( .INIT(8'h80) )  psh_negedge_reg_1_sqmuxa_8 (.A(
        PRDATA_regif_sn_m21_a0_0_net_1), .B(
        psh_negedge_reg_1_sqmuxa_8_1_0), .C(psh_prescale_reg13_net_1), 
        .Y(psh_negedge_reg_1_sqmuxa_8_net_1));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[13]  (.A(
        pwm_negedge_reg[142]), .B(pwm_negedge_reg[94]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_741));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_12  (.A(period_reg[12])
        , .B(period_cnt[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_11), .S(), .Y(), .FCO(un1_period_cnt_cry_12)
        );
    CFG2 #( .INIT(4'h8) )  psh_negedge_reg_1_sqmuxa_2_2 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        psh_negedge_reg_1_sqmuxa_3_2));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_1[2]  (.A(
        pwm_negedge_reg[83]), .B(pwm_enable_reg[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\PRDATA_regif_12_1_0[2] ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[33]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[33]));
    CFG4 #( .INIT(16'h1903) )  PRDATA_regif_sn_m25_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        PRDATA_regif_sn_m25_1_net_1));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[55]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[55]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[41]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[41]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[19]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[19]));
    CFG4 #( .INIT(16'h93C7) )  PRDATA_regif_sn_m25 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        PRDATA_regif_sn_m25_1_net_1), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(PRDATA_regif_sn_N_26));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[13]  (.A(
        pwm_negedge_reg[158]), .B(pwm_negedge_reg[30]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[13]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[11]  (.A(N_775), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_791), .Y(N_829));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[49]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[49]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[110]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[110]));
    CFG3 #( .INIT(8'h80) )  psh_negedge_reg_1_sqmuxa_6 (.A(
        PRDATA_regif_sn_m21_a0_0_net_1), .B(
        psh_negedge_reg_1_sqmuxa_6_1_net_1), .C(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_6_net_1)
        );
    SLE \psh_enable_reg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[7]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[122]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[122]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_0[1]  (.A(
        pwm_negedge_reg[130]), .B(period_reg[1]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\PRDATA_regif_12_1[1] ));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[3]  (.A(
        pwm_negedge_reg[36]), .B(pwm_negedge_reg[100]), .C(
        \PRDATA_regif_10_1_1[3] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_767));
    CFG4 #( .INIT(16'h0040) )  psh_negedge_reg_1_sqmuxa_1_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        psh_negedge_reg_1_sqmuxa_1_0_net_1));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[15]  (.A(
        pwm_negedge_reg[144]), .B(pwm_negedge_reg[96]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_743));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[8]  (.A(N_736), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[8]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_806));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[15]  (.A(
        pwm_negedge_reg[48]), .B(pwm_negedge_reg[112]), .C(
        \PRDATA_regif_10_1_1[15] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_779));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[81]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[81]));
    SLE \psh_period_reg[9]  (.D(CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[9]_net_1 ));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[15]  (.A(N_743), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[15]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_813));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[130]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[130]));
    CFG3 #( .INIT(8'h10) )  \PRDATA_regif_9[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[7]), .B(un1_OEn_2), .C(
        \PRDATA_regif_9_1[0]_net_1 ), .Y(N_762));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[4]  (.A(N_768), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_784), .Y(N_822));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[14]  (.A(
        pwm_negedge_reg[63]), .B(pwm_negedge_reg[127]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[14] ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_15_bm[5]  (.A(N_769), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_785), .Y(
        \PRDATA_regif_15_bm[5]_net_1 ));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[15]  (.A(
        pwm_negedge_reg[64]), .B(pwm_negedge_reg[128]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[15] ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[39]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[39]));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_am_1[5]  (.A(
        pwm_negedge_reg[134]), .B(period_reg[5]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_15_am_1[5]_net_1 ));
    SLE \period_reg[1]  (.D(\psh_period_reg[1]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[1]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[66]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[66]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_13  (.A(period_reg[13])
        , .B(period_cnt[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_12), .S(), .Y(), .FCO(un1_period_cnt_cry_13)
        );
    SLE \period_reg[6]  (.D(\psh_period_reg[6]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[6]));
    SLE \psh_enable_reg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[1]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[30]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[30]));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_RNO[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\PRDATA_regif_12_1[3] ), 
        .C(\PRDATA_regif_12_1_0[3] ), .Y(N_801));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[9]  (.A(
        \PRDATA_regif_11_bm[9]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[9]_net_1 ), .Y(N_789));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[9]  (.A(N_737), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[9]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_807));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[7]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[7]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[145]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[145]));
    CFG3 #( .INIT(8'h40) )  psh_negedge_reg_1_sqmuxa_1 (.A(
        un3_PRDATA_regif_1), .B(psh_negedge_reg_1_sqmuxa_1_0_net_1), 
        .C(psh_prescale_reg13_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'h7000) )  \PRDATA_regif_9_1[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(pwm_enable_reg[9]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_regif_9_1[0]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[76]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[76]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[17]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[17]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[156]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[156]));
    CFG4 #( .INIT(16'h1000) )  psh_enable_reg2_1_sqmuxa (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_enable_reg2_1_sqmuxa_1_0_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_enable_reg2_1_sqmuxa_net_1));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[53]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[53]));
    SLE \psh_enable_reg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[5]));
    SLE \psh_enable_reg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[3]));
    SLE \psh_enable_reg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[2]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[100]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[100]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[54]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[54]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_0  (.A(period_reg[0]), 
        .B(period_cnt[0]), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(un1_period_cnt_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_9  (.A(period_reg[9]), 
        .B(period_cnt[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_8), .S(), .Y(), .FCO(un1_period_cnt_cry_9));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[83]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[83]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[91]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[91]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[124]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[124]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[140]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[140]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[160]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[160]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[6]  (.A(
        pwm_negedge_reg[71]), .B(pwm_negedge_reg[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[6]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[12]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[12]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[15]  (.A(
        pwm_negedge_reg[160]), .B(pwm_negedge_reg[32]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[15]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[61]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[61]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[10]  (.A(
        pwm_negedge_reg[59]), .B(pwm_negedge_reg[123]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[10] ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[112]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[112]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_am[3]  (.A(
        pwm_negedge_reg[68]), .B(pwm_negedge_reg[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        \PRDATA_regif_11_am[3]_net_1 ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[90]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[90]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[128]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[128]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[158]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[158]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[117]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[117]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[132]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[132]));
    CFG3 #( .INIT(8'h80) )  psh_negedge_reg_1_sqmuxa_8_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        psh_negedge_reg_1_sqmuxa_8_1_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_8_1_0));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[3]  (.A(
        \PRDATA_regif_11_bm[3]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[3]_net_1 ), .Y(N_783));
    SLE \psh_period_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[3]_net_1 ));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_1[0]  (.A(
        pwm_negedge_reg[81]), .B(pwm_enable_reg[1]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\PRDATA_regif_12_1_0[0] ));
    CFG3 #( .INIT(8'h53) )  \PRDATA_regif_15_RNO_0[2]  (.A(
        pwm_negedge_reg[131]), .B(period_reg[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(\PRDATA_regif_12_1[2] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_10  (.A(period_reg[10])
        , .B(period_cnt[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_9), .S(), .Y(), .FCO(un1_period_cnt_cry_10));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[13]  (.A(
        pwm_negedge_reg[62]), .B(pwm_negedge_reg[126]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[13] ));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[12]  (.A(
        pwm_negedge_reg[141]), .B(pwm_negedge_reg[93]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_740));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[139]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[139]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[93]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[93]));
    SLE \psh_period_reg[15]  (.D(CoreAPB3_0_APBmslave0_PWDATA[15]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[15]_net_1 )
        );
    CFG4 #( .INIT(16'h0010) )  psh_period_reg_1_sqmuxa_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        psh_period_reg_1_sqmuxa_1_net_1));
    CFG2 #( .INIT(4'h4) )  psh_negedge_reg_1_sqmuxa_2_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        psh_negedge_reg_1_sqmuxa_8_1_net_1));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[11]  (.A(
        pwm_negedge_reg[156]), .B(pwm_negedge_reg[28]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[11]_net_1 ));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[4]  (.A(
        pwm_negedge_reg[53]), .B(pwm_negedge_reg[117]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[4] ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[102]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[102]));
    CFG4 #( .INIT(16'h4000) )  psh_negedge_reg_1_sqmuxa_5 (.A(
        un3_PRDATA_regif_1), .B(psh_negedge_reg_1_sqmuxa_5_2), .C(
        psh_prescale_reg13_net_1), .D(
        psh_negedge_reg_1_sqmuxa_8_1_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_5_net_1));
    CFG3 #( .INIT(8'h80) )  psh_negedge_reg_1_sqmuxa_4_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        psh_negedge_reg_1_sqmuxa_8_1_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_4_1_net_1));
    CFG4 #( .INIT(16'h0008) )  psh_enable_reg2_1_sqmuxa_1_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        psh_enable_reg2_1_sqmuxa_1_0_net_1));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[86]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[86]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_15_bm_RNO_0[5]  (.A(
        pwm_negedge_reg[54]), .B(pwm_negedge_reg[118]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[5] ));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[0]  (.A(
        pwm_negedge_reg[49]), .B(pwm_negedge_reg[113]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1[0] ));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[142]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[142]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[1]  (.A(
        \PRDATA_regif_11_bm[1]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[1]_net_1 ), .Y(N_781));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[10]  (.A(
        \PRDATA_regif_11_bm[10]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[10]_net_1 ), .Y(N_790));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[21]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[21]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[113]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[113]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[109]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[109]));
    CFG4 #( .INIT(16'h8000) )  psh_prescale_reg13 (.A(
        CoreAPB3_0_APBmslave0_PENABLE), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .C(iPSELS_0_0[4]), .D(
        iPSELS_0[4]), .Y(psh_prescale_reg13_net_1));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[134]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[134]));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_RNO[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\PRDATA_regif_12_1[1] ), 
        .C(\PRDATA_regif_12_1_0[1] ), .Y(N_799));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[9]  (.A(
        pwm_negedge_reg[154]), .B(pwm_negedge_reg[26]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[9]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[14]  (.A(N_778), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_794), .Y(N_832));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[146]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[146]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[5]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[5]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[16]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[16]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[10]  (.A(N_774), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_790), .Y(N_828));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[72]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[72]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[48]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[48]));
    CFG4 #( .INIT(16'hEFFF) )  PRDATA_regif_13_N_5L8 (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(controlReg14_3), .D(
        PRDATA_regif_sn_m21_a0_0_net_1), .Y(
        PRDATA_regif_13_N_5L8_net_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_6  (.A(period_reg[6]), 
        .B(period_cnt[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_5), .S(), .Y(), .FCO(un1_period_cnt_cry_6));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[138]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[138]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[98]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[98]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[24]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[24]));
    SLE \psh_period_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[4]_net_1 ));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[8]  (.A(
        pwm_negedge_reg[41]), .B(pwm_negedge_reg[105]), .C(
        \PRDATA_regif_10_1_1[8] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_772));
    CFG4 #( .INIT(16'h0FCA) )  \PRDATA_regif_14_RNO[9]  (.A(
        pwm_negedge_reg[42]), .B(pwm_negedge_reg[106]), .C(
        \PRDATA_regif_10_1_1[9] ), .D(CoreAPB3_0_APBmslave0_PADDR[3]), 
        .Y(N_773));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[152]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[152]));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[11]  (.A(
        pwm_negedge_reg[60]), .B(pwm_negedge_reg[124]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[11] ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[96]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[96]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[104]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[104]));
    CFG3 #( .INIT(8'hCA) )  \PRDATA_regif_7[11]  (.A(
        pwm_negedge_reg[140]), .B(pwm_negedge_reg[92]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_739));
    CFG4 #( .INIT(16'h8000) )  psh_negedge_reg_1_sqmuxa_2 (.A(
        psh_negedge_reg_1_sqmuxa_3_2), .B(psh_negedge_reg_1_sqmuxa_5_2)
        , .C(psh_prescale_reg13_net_1), .D(
        psh_negedge_reg_1_sqmuxa_8_1_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_2_net_1));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[32]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[32]));
    CFG3 #( .INIT(8'h80) )  psh_negedge_reg_1_sqmuxa_7 (.A(
        PRDATA_regif_sn_m21_a0_0_net_1), .B(
        psh_negedge_reg_1_sqmuxa_7_1_net_1), .C(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_7_net_1)
        );
    SLE \period_reg[7]  (.D(\psh_period_reg[7]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[7]));
    SLE \psh_period_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[7]_net_1 ));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_RNO[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\PRDATA_regif_12_1[2] ), 
        .C(\PRDATA_regif_12_1_0[2] ), .Y(N_800));
    CFG4 #( .INIT(16'h530F) )  \PRDATA_regif_14_RNO_0[9]  (.A(
        pwm_negedge_reg[58]), .B(pwm_negedge_reg[122]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_10_1_1[9] ));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_14[13]  (.A(N_777), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_793), .Y(N_831));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[144]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[144]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[148]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[148]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[108]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[108]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[74]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[74]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[0]  (.A(
        pwm_negedge_reg[145]), .B(pwm_negedge_reg[17]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[0]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[51]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[51]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[67]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[67]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[56]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[56]));
    SLE \period_reg[10]  (.D(\psh_period_reg[10]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[10]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[121]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[121]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_15_bm[7]  (.A(N_771), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(N_787), .Y(
        \PRDATA_regif_15_bm[7]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[77]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_8_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[77]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[26]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[26]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[5]  (.A(
        pwm_negedge_reg[150]), .B(pwm_negedge_reg[22]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[5]_net_1 ));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[29]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[29]));
    SLE \psh_enable_reg2[10]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), 
        .CLK(GL0_INST), .EN(psh_enable_reg2_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[10]));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_RNO[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\PRDATA_regif_12_1[0] ), 
        .C(\PRDATA_regif_12_1_0[0] ), .Y(N_798));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[59]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[59]));
    SLE \psh_enable_reg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[6]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[6]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[6]));
    CFG3 #( .INIT(8'h1B) )  \PRDATA_regif_15_am[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        \PRDATA_regif_15_am_1[5]_net_1 ), .C(
        \PRDATA_regif_15_am_1_0[5]_net_1 ), .Y(
        \PRDATA_regif_15_am[5]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[14]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[14]));
    SLE \gen_pos_neg_shregs[9].psh_negedge_reg[129]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[129]));
    CFG4 #( .INIT(16'h292A) )  PRDATA_regif_sn_m31 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .D(controlReg24_3), .Y(
        PRDATA_regif_sn_N_39_mux));
    CFG3 #( .INIT(8'h40) )  psh_period_reg_1_sqmuxa (.A(
        un3_PRDATA_regif_1), .B(psh_period_reg_1_sqmuxa_1_net_1), .C(
        psh_prescale_reg13_net_1), .Y(psh_period_reg_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'h0004) )  psh_enable_reg1_1_sqmuxa_2 (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        CoreAPB3_0_APBmslave0_PADDR[5]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        psh_enable_reg1_1_sqmuxa_2_net_1));
    SLE \psh_enable_reg2[9]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), 
        .CLK(GL0_INST), .EN(psh_enable_reg2_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[9]));
    SLE \psh_period_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[6]_net_1 ));
    CFG4 #( .INIT(16'h22E2) )  \PRDATA_regif_12[11]  (.A(N_739), .B(
        PRDATA_regif_sn_N_15), .C(period_reg[11]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_809));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[18]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_9_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[18]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[2]  (.A(
        \PRDATA_regif_11_bm[2]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        \PRDATA_regif_11_am[2]_net_1 ), .Y(N_782));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[47]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[47]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[125]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[125]));
    SLE \period_reg[15]  (.D(\psh_period_reg[15]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[15]));
    SLE \gen_pos_neg_shregs[10].psh_negedge_reg[159]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[159]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[38]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[38]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_11_bm[4]  (.A(
        pwm_negedge_reg[149]), .B(pwm_negedge_reg[21]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(
        \PRDATA_regif_11_bm[4]_net_1 ));
    
endmodule


module corepwm_Z5(
       CoreAPB3_0_APBmslave0_PWDATA,
       iPSELS_0_0,
       iPSELS_0,
       CoreAPB3_0_APBmslave0_PADDR,
       CoreAPB3_0_APBmslave4_PRDATA,
       PWM_c,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       N_97_1,
       controlReg14_3,
       PRDATA_regif_sn_N_26,
       N_842,
       N_841,
       N_840,
       un1_OEn_2,
       un3_PRDATA_regif_1,
       psh_negedge_reg_1_sqmuxa_3_2,
       N_813,
       N_811,
       N_806,
       N_812,
       N_807,
       N_808,
       N_810,
       N_809,
       controlReg24_3,
       PRDATA_regif_sn_N_39_mux,
       N_833,
       N_831,
       N_828,
       N_826,
       N_832,
       N_827,
       N_830,
       N_829,
       N_837,
       N_839,
       N_838
    );
input  [15:0] CoreAPB3_0_APBmslave0_PWDATA;
input  [4:4] iPSELS_0_0;
input  [4:4] iPSELS_0;
input  [7:2] CoreAPB3_0_APBmslave0_PADDR;
output [1:0] CoreAPB3_0_APBmslave4_PRDATA;
output [10:1] PWM_c;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  N_97_1;
input  controlReg14_3;
output PRDATA_regif_sn_N_26;
output N_842;
output N_841;
output N_840;
input  un1_OEn_2;
output un3_PRDATA_regif_1;
output psh_negedge_reg_1_sqmuxa_3_2;
output N_813;
output N_811;
output N_806;
output N_812;
output N_807;
output N_808;
output N_810;
output N_809;
input  controlReg24_3;
output PRDATA_regif_sn_N_39_mux;
output N_833;
output N_831;
output N_828;
output N_826;
output N_832;
output N_827;
output N_830;
output N_829;
output N_837;
output N_839;
output N_838;

    wire \pwm_enable_reg[1] , \pwm_enable_reg[2] , \pwm_enable_reg[3] , 
        \pwm_enable_reg[4] , \pwm_enable_reg[5] , \pwm_enable_reg[6] , 
        \pwm_enable_reg[7] , \pwm_enable_reg[8] , \pwm_enable_reg[9] , 
        \pwm_enable_reg[10] , \pwm_negedge_reg[1] , 
        \pwm_negedge_reg[2] , \pwm_negedge_reg[3] , 
        \pwm_negedge_reg[4] , \pwm_negedge_reg[5] , 
        \pwm_negedge_reg[6] , \pwm_negedge_reg[7] , 
        \pwm_negedge_reg[8] , \pwm_negedge_reg[9] , 
        \pwm_negedge_reg[10] , \pwm_negedge_reg[11] , 
        \pwm_negedge_reg[12] , \pwm_negedge_reg[13] , 
        \pwm_negedge_reg[14] , \pwm_negedge_reg[15] , 
        \pwm_negedge_reg[16] , \pwm_negedge_reg[17] , 
        \pwm_negedge_reg[18] , \pwm_negedge_reg[19] , 
        \pwm_negedge_reg[20] , \pwm_negedge_reg[21] , 
        \pwm_negedge_reg[22] , \pwm_negedge_reg[23] , 
        \pwm_negedge_reg[24] , \pwm_negedge_reg[25] , 
        \pwm_negedge_reg[26] , \pwm_negedge_reg[27] , 
        \pwm_negedge_reg[28] , \pwm_negedge_reg[29] , 
        \pwm_negedge_reg[30] , \pwm_negedge_reg[31] , 
        \pwm_negedge_reg[32] , \pwm_negedge_reg[33] , 
        \pwm_negedge_reg[34] , \pwm_negedge_reg[35] , 
        \pwm_negedge_reg[36] , \pwm_negedge_reg[37] , 
        \pwm_negedge_reg[38] , \pwm_negedge_reg[39] , 
        \pwm_negedge_reg[40] , \pwm_negedge_reg[41] , 
        \pwm_negedge_reg[42] , \pwm_negedge_reg[43] , 
        \pwm_negedge_reg[44] , \pwm_negedge_reg[45] , 
        \pwm_negedge_reg[46] , \pwm_negedge_reg[47] , 
        \pwm_negedge_reg[48] , \pwm_negedge_reg[49] , 
        \pwm_negedge_reg[50] , \pwm_negedge_reg[51] , 
        \pwm_negedge_reg[52] , \pwm_negedge_reg[53] , 
        \pwm_negedge_reg[54] , \pwm_negedge_reg[55] , 
        \pwm_negedge_reg[56] , \pwm_negedge_reg[57] , 
        \pwm_negedge_reg[58] , \pwm_negedge_reg[59] , 
        \pwm_negedge_reg[60] , \pwm_negedge_reg[61] , 
        \pwm_negedge_reg[62] , \pwm_negedge_reg[63] , 
        \pwm_negedge_reg[64] , \pwm_negedge_reg[65] , 
        \pwm_negedge_reg[66] , \pwm_negedge_reg[67] , 
        \pwm_negedge_reg[68] , \pwm_negedge_reg[69] , 
        \pwm_negedge_reg[70] , \pwm_negedge_reg[71] , 
        \pwm_negedge_reg[72] , \pwm_negedge_reg[73] , 
        \pwm_negedge_reg[74] , \pwm_negedge_reg[75] , 
        \pwm_negedge_reg[76] , \pwm_negedge_reg[77] , 
        \pwm_negedge_reg[78] , \pwm_negedge_reg[79] , 
        \pwm_negedge_reg[80] , \pwm_negedge_reg[81] , 
        \pwm_negedge_reg[82] , \pwm_negedge_reg[83] , 
        \pwm_negedge_reg[84] , \pwm_negedge_reg[85] , 
        \pwm_negedge_reg[86] , \pwm_negedge_reg[87] , 
        \pwm_negedge_reg[88] , \pwm_negedge_reg[89] , 
        \pwm_negedge_reg[90] , \pwm_negedge_reg[91] , 
        \pwm_negedge_reg[92] , \pwm_negedge_reg[93] , 
        \pwm_negedge_reg[94] , \pwm_negedge_reg[95] , 
        \pwm_negedge_reg[96] , \pwm_negedge_reg[97] , 
        \pwm_negedge_reg[98] , \pwm_negedge_reg[99] , 
        \pwm_negedge_reg[100] , \pwm_negedge_reg[101] , 
        \pwm_negedge_reg[102] , \pwm_negedge_reg[103] , 
        \pwm_negedge_reg[104] , \pwm_negedge_reg[105] , 
        \pwm_negedge_reg[106] , \pwm_negedge_reg[107] , 
        \pwm_negedge_reg[108] , \pwm_negedge_reg[109] , 
        \pwm_negedge_reg[110] , \pwm_negedge_reg[111] , 
        \pwm_negedge_reg[112] , \pwm_negedge_reg[113] , 
        \pwm_negedge_reg[114] , \pwm_negedge_reg[115] , 
        \pwm_negedge_reg[116] , \pwm_negedge_reg[117] , 
        \pwm_negedge_reg[118] , \pwm_negedge_reg[119] , 
        \pwm_negedge_reg[120] , \pwm_negedge_reg[121] , 
        \pwm_negedge_reg[122] , \pwm_negedge_reg[123] , 
        \pwm_negedge_reg[124] , \pwm_negedge_reg[125] , 
        \pwm_negedge_reg[126] , \pwm_negedge_reg[127] , 
        \pwm_negedge_reg[128] , \pwm_negedge_reg[129] , 
        \pwm_negedge_reg[130] , \pwm_negedge_reg[131] , 
        \pwm_negedge_reg[132] , \pwm_negedge_reg[133] , 
        \pwm_negedge_reg[134] , \pwm_negedge_reg[135] , 
        \pwm_negedge_reg[136] , \pwm_negedge_reg[137] , 
        \pwm_negedge_reg[138] , \pwm_negedge_reg[139] , 
        \pwm_negedge_reg[140] , \pwm_negedge_reg[141] , 
        \pwm_negedge_reg[142] , \pwm_negedge_reg[143] , 
        \pwm_negedge_reg[144] , \pwm_negedge_reg[145] , 
        \pwm_negedge_reg[146] , \pwm_negedge_reg[147] , 
        \pwm_negedge_reg[148] , \pwm_negedge_reg[149] , 
        \pwm_negedge_reg[150] , \pwm_negedge_reg[151] , 
        \pwm_negedge_reg[152] , \pwm_negedge_reg[153] , 
        \pwm_negedge_reg[154] , \pwm_negedge_reg[155] , 
        \pwm_negedge_reg[156] , \pwm_negedge_reg[157] , 
        \pwm_negedge_reg[158] , \pwm_negedge_reg[159] , 
        \pwm_negedge_reg[160] , \period_reg[0] , \period_reg[1] , 
        \period_reg[2] , \period_reg[3] , \period_reg[4] , 
        \period_reg[5] , \period_reg[6] , \period_reg[7] , 
        \period_reg[8] , \period_reg[9] , \period_reg[10] , 
        \period_reg[11] , \period_reg[12] , \period_reg[13] , 
        \period_reg[14] , \period_reg[15] , \period_cnt[0] , 
        \period_cnt[1] , \period_cnt[2] , \period_cnt[3] , 
        \period_cnt[4] , \period_cnt[5] , \period_cnt[6] , 
        \period_cnt[7] , \period_cnt[8] , \period_cnt[9] , 
        \period_cnt[10] , \period_cnt[11] , \period_cnt[12] , 
        \period_cnt[13] , \period_cnt[14] , \period_cnt[15] , 
        GND_net_1, VCC_net_1;
    
    pwm_gen_10s_16s_0 \genblk5.pwm_gen  (.PWM_c({PWM_c[10], PWM_c[9], 
        PWM_c[8], PWM_c[7], PWM_c[6], PWM_c[5], PWM_c[4], PWM_c[3], 
        PWM_c[2], PWM_c[1]}), .period_cnt({\period_cnt[15] , 
        \period_cnt[14] , \period_cnt[13] , \period_cnt[12] , 
        \period_cnt[11] , \period_cnt[10] , \period_cnt[9] , 
        \period_cnt[8] , \period_cnt[7] , \period_cnt[6] , 
        \period_cnt[5] , \period_cnt[4] , \period_cnt[3] , 
        \period_cnt[2] , \period_cnt[1] , \period_cnt[0] }), 
        .pwm_negedge_reg({\pwm_negedge_reg[160] , 
        \pwm_negedge_reg[159] , \pwm_negedge_reg[158] , 
        \pwm_negedge_reg[157] , \pwm_negedge_reg[156] , 
        \pwm_negedge_reg[155] , \pwm_negedge_reg[154] , 
        \pwm_negedge_reg[153] , \pwm_negedge_reg[152] , 
        \pwm_negedge_reg[151] , \pwm_negedge_reg[150] , 
        \pwm_negedge_reg[149] , \pwm_negedge_reg[148] , 
        \pwm_negedge_reg[147] , \pwm_negedge_reg[146] , 
        \pwm_negedge_reg[145] , \pwm_negedge_reg[144] , 
        \pwm_negedge_reg[143] , \pwm_negedge_reg[142] , 
        \pwm_negedge_reg[141] , \pwm_negedge_reg[140] , 
        \pwm_negedge_reg[139] , \pwm_negedge_reg[138] , 
        \pwm_negedge_reg[137] , \pwm_negedge_reg[136] , 
        \pwm_negedge_reg[135] , \pwm_negedge_reg[134] , 
        \pwm_negedge_reg[133] , \pwm_negedge_reg[132] , 
        \pwm_negedge_reg[131] , \pwm_negedge_reg[130] , 
        \pwm_negedge_reg[129] , \pwm_negedge_reg[128] , 
        \pwm_negedge_reg[127] , \pwm_negedge_reg[126] , 
        \pwm_negedge_reg[125] , \pwm_negedge_reg[124] , 
        \pwm_negedge_reg[123] , \pwm_negedge_reg[122] , 
        \pwm_negedge_reg[121] , \pwm_negedge_reg[120] , 
        \pwm_negedge_reg[119] , \pwm_negedge_reg[118] , 
        \pwm_negedge_reg[117] , \pwm_negedge_reg[116] , 
        \pwm_negedge_reg[115] , \pwm_negedge_reg[114] , 
        \pwm_negedge_reg[113] , \pwm_negedge_reg[112] , 
        \pwm_negedge_reg[111] , \pwm_negedge_reg[110] , 
        \pwm_negedge_reg[109] , \pwm_negedge_reg[108] , 
        \pwm_negedge_reg[107] , \pwm_negedge_reg[106] , 
        \pwm_negedge_reg[105] , \pwm_negedge_reg[104] , 
        \pwm_negedge_reg[103] , \pwm_negedge_reg[102] , 
        \pwm_negedge_reg[101] , \pwm_negedge_reg[100] , 
        \pwm_negedge_reg[99] , \pwm_negedge_reg[98] , 
        \pwm_negedge_reg[97] , \pwm_negedge_reg[96] , 
        \pwm_negedge_reg[95] , \pwm_negedge_reg[94] , 
        \pwm_negedge_reg[93] , \pwm_negedge_reg[92] , 
        \pwm_negedge_reg[91] , \pwm_negedge_reg[90] , 
        \pwm_negedge_reg[89] , \pwm_negedge_reg[88] , 
        \pwm_negedge_reg[87] , \pwm_negedge_reg[86] , 
        \pwm_negedge_reg[85] , \pwm_negedge_reg[84] , 
        \pwm_negedge_reg[83] , \pwm_negedge_reg[82] , 
        \pwm_negedge_reg[81] , \pwm_negedge_reg[80] , 
        \pwm_negedge_reg[79] , \pwm_negedge_reg[78] , 
        \pwm_negedge_reg[77] , \pwm_negedge_reg[76] , 
        \pwm_negedge_reg[75] , \pwm_negedge_reg[74] , 
        \pwm_negedge_reg[73] , \pwm_negedge_reg[72] , 
        \pwm_negedge_reg[71] , \pwm_negedge_reg[70] , 
        \pwm_negedge_reg[69] , \pwm_negedge_reg[68] , 
        \pwm_negedge_reg[67] , \pwm_negedge_reg[66] , 
        \pwm_negedge_reg[65] , \pwm_negedge_reg[64] , 
        \pwm_negedge_reg[63] , \pwm_negedge_reg[62] , 
        \pwm_negedge_reg[61] , \pwm_negedge_reg[60] , 
        \pwm_negedge_reg[59] , \pwm_negedge_reg[58] , 
        \pwm_negedge_reg[57] , \pwm_negedge_reg[56] , 
        \pwm_negedge_reg[55] , \pwm_negedge_reg[54] , 
        \pwm_negedge_reg[53] , \pwm_negedge_reg[52] , 
        \pwm_negedge_reg[51] , \pwm_negedge_reg[50] , 
        \pwm_negedge_reg[49] , \pwm_negedge_reg[48] , 
        \pwm_negedge_reg[47] , \pwm_negedge_reg[46] , 
        \pwm_negedge_reg[45] , \pwm_negedge_reg[44] , 
        \pwm_negedge_reg[43] , \pwm_negedge_reg[42] , 
        \pwm_negedge_reg[41] , \pwm_negedge_reg[40] , 
        \pwm_negedge_reg[39] , \pwm_negedge_reg[38] , 
        \pwm_negedge_reg[37] , \pwm_negedge_reg[36] , 
        \pwm_negedge_reg[35] , \pwm_negedge_reg[34] , 
        \pwm_negedge_reg[33] , \pwm_negedge_reg[32] , 
        \pwm_negedge_reg[31] , \pwm_negedge_reg[30] , 
        \pwm_negedge_reg[29] , \pwm_negedge_reg[28] , 
        \pwm_negedge_reg[27] , \pwm_negedge_reg[26] , 
        \pwm_negedge_reg[25] , \pwm_negedge_reg[24] , 
        \pwm_negedge_reg[23] , \pwm_negedge_reg[22] , 
        \pwm_negedge_reg[21] , \pwm_negedge_reg[20] , 
        \pwm_negedge_reg[19] , \pwm_negedge_reg[18] , 
        \pwm_negedge_reg[17] , \pwm_negedge_reg[16] , 
        \pwm_negedge_reg[15] , \pwm_negedge_reg[14] , 
        \pwm_negedge_reg[13] , \pwm_negedge_reg[12] , 
        \pwm_negedge_reg[11] , \pwm_negedge_reg[10] , 
        \pwm_negedge_reg[9] , \pwm_negedge_reg[8] , 
        \pwm_negedge_reg[7] , \pwm_negedge_reg[6] , 
        \pwm_negedge_reg[5] , \pwm_negedge_reg[4] , 
        \pwm_negedge_reg[3] , \pwm_negedge_reg[2] , 
        \pwm_negedge_reg[1] }), .pwm_enable_reg({\pwm_enable_reg[10] , 
        \pwm_enable_reg[9] , \pwm_enable_reg[8] , \pwm_enable_reg[7] , 
        \pwm_enable_reg[6] , \pwm_enable_reg[5] , \pwm_enable_reg[4] , 
        \pwm_enable_reg[3] , \pwm_enable_reg[2] , \pwm_enable_reg[1] })
        , .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    timebase_16s \genblk4.genblk1.timebase  (.period_cnt({
        \period_cnt[15] , \period_cnt[14] , \period_cnt[13] , 
        \period_cnt[12] , \period_cnt[11] , \period_cnt[10] , 
        \period_cnt[9] , \period_cnt[8] , \period_cnt[7] , 
        \period_cnt[6] , \period_cnt[5] , \period_cnt[4] , 
        \period_cnt[3] , \period_cnt[2] , \period_cnt[1] , 
        \period_cnt[0] }), .period_reg({\period_reg[15] , 
        \period_reg[14] , \period_reg[13] , \period_reg[12] , 
        \period_reg[11] , \period_reg[10] , \period_reg[9] , 
        \period_reg[8] , \period_reg[7] , \period_reg[6] , 
        \period_reg[5] , \period_reg[4] , \period_reg[3] , 
        \period_reg[2] , \period_reg[1] , \period_reg[0] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST));
    reg_if_Z6 \genblk2.reg_if  (.CoreAPB3_0_APBmslave0_PWDATA({
        CoreAPB3_0_APBmslave0_PWDATA[15], 
        CoreAPB3_0_APBmslave0_PWDATA[14], 
        CoreAPB3_0_APBmslave0_PWDATA[13], 
        CoreAPB3_0_APBmslave0_PWDATA[12], 
        CoreAPB3_0_APBmslave0_PWDATA[11], 
        CoreAPB3_0_APBmslave0_PWDATA[10], 
        CoreAPB3_0_APBmslave0_PWDATA[9], 
        CoreAPB3_0_APBmslave0_PWDATA[8], 
        CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .pwm_enable_reg({
        \pwm_enable_reg[10] , \pwm_enable_reg[9] , \pwm_enable_reg[8] , 
        \pwm_enable_reg[7] , \pwm_enable_reg[6] , \pwm_enable_reg[5] , 
        \pwm_enable_reg[4] , \pwm_enable_reg[3] , \pwm_enable_reg[2] , 
        \pwm_enable_reg[1] }), .pwm_negedge_reg({
        \pwm_negedge_reg[160] , \pwm_negedge_reg[159] , 
        \pwm_negedge_reg[158] , \pwm_negedge_reg[157] , 
        \pwm_negedge_reg[156] , \pwm_negedge_reg[155] , 
        \pwm_negedge_reg[154] , \pwm_negedge_reg[153] , 
        \pwm_negedge_reg[152] , \pwm_negedge_reg[151] , 
        \pwm_negedge_reg[150] , \pwm_negedge_reg[149] , 
        \pwm_negedge_reg[148] , \pwm_negedge_reg[147] , 
        \pwm_negedge_reg[146] , \pwm_negedge_reg[145] , 
        \pwm_negedge_reg[144] , \pwm_negedge_reg[143] , 
        \pwm_negedge_reg[142] , \pwm_negedge_reg[141] , 
        \pwm_negedge_reg[140] , \pwm_negedge_reg[139] , 
        \pwm_negedge_reg[138] , \pwm_negedge_reg[137] , 
        \pwm_negedge_reg[136] , \pwm_negedge_reg[135] , 
        \pwm_negedge_reg[134] , \pwm_negedge_reg[133] , 
        \pwm_negedge_reg[132] , \pwm_negedge_reg[131] , 
        \pwm_negedge_reg[130] , \pwm_negedge_reg[129] , 
        \pwm_negedge_reg[128] , \pwm_negedge_reg[127] , 
        \pwm_negedge_reg[126] , \pwm_negedge_reg[125] , 
        \pwm_negedge_reg[124] , \pwm_negedge_reg[123] , 
        \pwm_negedge_reg[122] , \pwm_negedge_reg[121] , 
        \pwm_negedge_reg[120] , \pwm_negedge_reg[119] , 
        \pwm_negedge_reg[118] , \pwm_negedge_reg[117] , 
        \pwm_negedge_reg[116] , \pwm_negedge_reg[115] , 
        \pwm_negedge_reg[114] , \pwm_negedge_reg[113] , 
        \pwm_negedge_reg[112] , \pwm_negedge_reg[111] , 
        \pwm_negedge_reg[110] , \pwm_negedge_reg[109] , 
        \pwm_negedge_reg[108] , \pwm_negedge_reg[107] , 
        \pwm_negedge_reg[106] , \pwm_negedge_reg[105] , 
        \pwm_negedge_reg[104] , \pwm_negedge_reg[103] , 
        \pwm_negedge_reg[102] , \pwm_negedge_reg[101] , 
        \pwm_negedge_reg[100] , \pwm_negedge_reg[99] , 
        \pwm_negedge_reg[98] , \pwm_negedge_reg[97] , 
        \pwm_negedge_reg[96] , \pwm_negedge_reg[95] , 
        \pwm_negedge_reg[94] , \pwm_negedge_reg[93] , 
        \pwm_negedge_reg[92] , \pwm_negedge_reg[91] , 
        \pwm_negedge_reg[90] , \pwm_negedge_reg[89] , 
        \pwm_negedge_reg[88] , \pwm_negedge_reg[87] , 
        \pwm_negedge_reg[86] , \pwm_negedge_reg[85] , 
        \pwm_negedge_reg[84] , \pwm_negedge_reg[83] , 
        \pwm_negedge_reg[82] , \pwm_negedge_reg[81] , 
        \pwm_negedge_reg[80] , \pwm_negedge_reg[79] , 
        \pwm_negedge_reg[78] , \pwm_negedge_reg[77] , 
        \pwm_negedge_reg[76] , \pwm_negedge_reg[75] , 
        \pwm_negedge_reg[74] , \pwm_negedge_reg[73] , 
        \pwm_negedge_reg[72] , \pwm_negedge_reg[71] , 
        \pwm_negedge_reg[70] , \pwm_negedge_reg[69] , 
        \pwm_negedge_reg[68] , \pwm_negedge_reg[67] , 
        \pwm_negedge_reg[66] , \pwm_negedge_reg[65] , 
        \pwm_negedge_reg[64] , \pwm_negedge_reg[63] , 
        \pwm_negedge_reg[62] , \pwm_negedge_reg[61] , 
        \pwm_negedge_reg[60] , \pwm_negedge_reg[59] , 
        \pwm_negedge_reg[58] , \pwm_negedge_reg[57] , 
        \pwm_negedge_reg[56] , \pwm_negedge_reg[55] , 
        \pwm_negedge_reg[54] , \pwm_negedge_reg[53] , 
        \pwm_negedge_reg[52] , \pwm_negedge_reg[51] , 
        \pwm_negedge_reg[50] , \pwm_negedge_reg[49] , 
        \pwm_negedge_reg[48] , \pwm_negedge_reg[47] , 
        \pwm_negedge_reg[46] , \pwm_negedge_reg[45] , 
        \pwm_negedge_reg[44] , \pwm_negedge_reg[43] , 
        \pwm_negedge_reg[42] , \pwm_negedge_reg[41] , 
        \pwm_negedge_reg[40] , \pwm_negedge_reg[39] , 
        \pwm_negedge_reg[38] , \pwm_negedge_reg[37] , 
        \pwm_negedge_reg[36] , \pwm_negedge_reg[35] , 
        \pwm_negedge_reg[34] , \pwm_negedge_reg[33] , 
        \pwm_negedge_reg[32] , \pwm_negedge_reg[31] , 
        \pwm_negedge_reg[30] , \pwm_negedge_reg[29] , 
        \pwm_negedge_reg[28] , \pwm_negedge_reg[27] , 
        \pwm_negedge_reg[26] , \pwm_negedge_reg[25] , 
        \pwm_negedge_reg[24] , \pwm_negedge_reg[23] , 
        \pwm_negedge_reg[22] , \pwm_negedge_reg[21] , 
        \pwm_negedge_reg[20] , \pwm_negedge_reg[19] , 
        \pwm_negedge_reg[18] , \pwm_negedge_reg[17] , 
        \pwm_negedge_reg[16] , \pwm_negedge_reg[15] , 
        \pwm_negedge_reg[14] , \pwm_negedge_reg[13] , 
        \pwm_negedge_reg[12] , \pwm_negedge_reg[11] , 
        \pwm_negedge_reg[10] , \pwm_negedge_reg[9] , 
        \pwm_negedge_reg[8] , \pwm_negedge_reg[7] , 
        \pwm_negedge_reg[6] , \pwm_negedge_reg[5] , 
        \pwm_negedge_reg[4] , \pwm_negedge_reg[3] , 
        \pwm_negedge_reg[2] , \pwm_negedge_reg[1] }), .period_reg({
        \period_reg[15] , \period_reg[14] , \period_reg[13] , 
        \period_reg[12] , \period_reg[11] , \period_reg[10] , 
        \period_reg[9] , \period_reg[8] , \period_reg[7] , 
        \period_reg[6] , \period_reg[5] , \period_reg[4] , 
        \period_reg[3] , \period_reg[2] , \period_reg[1] , 
        \period_reg[0] }), .period_cnt({\period_cnt[15] , 
        \period_cnt[14] , \period_cnt[13] , \period_cnt[12] , 
        \period_cnt[11] , \period_cnt[10] , \period_cnt[9] , 
        \period_cnt[8] , \period_cnt[7] , \period_cnt[6] , 
        \period_cnt[5] , \period_cnt[4] , \period_cnt[3] , 
        \period_cnt[2] , \period_cnt[1] , \period_cnt[0] }), 
        .iPSELS_0_0({iPSELS_0_0[4]}), .iPSELS_0({iPSELS_0[4]}), 
        .CoreAPB3_0_APBmslave0_PADDR({CoreAPB3_0_APBmslave0_PADDR[7], 
        CoreAPB3_0_APBmslave0_PADDR[6], CoreAPB3_0_APBmslave0_PADDR[5], 
        CoreAPB3_0_APBmslave0_PADDR[4], CoreAPB3_0_APBmslave0_PADDR[3], 
        CoreAPB3_0_APBmslave0_PADDR[2]}), 
        .CoreAPB3_0_APBmslave4_PRDATA({CoreAPB3_0_APBmslave4_PRDATA[1], 
        CoreAPB3_0_APBmslave4_PRDATA[0]}), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .N_97_1(N_97_1), .controlReg14_3(controlReg14_3), 
        .PRDATA_regif_sn_N_26(PRDATA_regif_sn_N_26), .N_842(N_842), 
        .N_841(N_841), .N_840(N_840), .un1_OEn_2(un1_OEn_2), 
        .un3_PRDATA_regif_1(un3_PRDATA_regif_1), 
        .psh_negedge_reg_1_sqmuxa_3_2(psh_negedge_reg_1_sqmuxa_3_2), 
        .N_813(N_813), .N_811(N_811), .N_806(N_806), .N_812(N_812), 
        .N_807(N_807), .N_808(N_808), .N_810(N_810), .N_809(N_809), 
        .controlReg24_3(controlReg24_3), .PRDATA_regif_sn_N_39_mux(
        PRDATA_regif_sn_N_39_mux), .N_833(N_833), .N_831(N_831), 
        .N_828(N_828), .N_826(N_826), .N_832(N_832), .N_827(N_827), 
        .N_830(N_830), .N_829(N_829), .N_837(N_837), .N_839(N_839), 
        .N_838(N_838));
    
endmodule


module mss_sb_MSS(
       CoreAPB3_0_APBmslave0_PADDR,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR,
       CoreAPB3_0_APBmslave0_PWDATA,
       COREI2C_0_0_INT,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N,
       CoreAPB3_0_APBmslave0_PENABLE,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       mss_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       CoreUARTapb_2_0_intr_or_2_Y,
       CoreUARTapb_2_1_intr_or_2_Y,
       LOCK,
       GL0_INST
    );
output [8:0] CoreAPB3_0_APBmslave0_PADDR;
output [15:12] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR;
output [15:0] CoreAPB3_0_APBmslave0_PWDATA;
input  [0:0] COREI2C_0_0_INT;
input  [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
output mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N;
output CoreAPB3_0_APBmslave0_PENABLE;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave0_PWRITE;
output mss_sb_MSS_TMP_0_MSS_RESET_N_M2F;
input  CoreUARTapb_2_0_intr_or_2_Y;
input  CoreUARTapb_2_1_intr_or_2_Y;
input  LOCK;
input  GL0_INST;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    MSS_010 #( .INIT(1438'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C00000000609300000003FFFFE400000000000010000000000F01C000001FEDFFC010842108421000001FE34001FF8000000400000000020051007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(0.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, 
        nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12], nc56, nc57, nc58, 
        CoreAPB3_0_APBmslave0_PADDR[8], CoreAPB3_0_APBmslave0_PADDR[7], 
        CoreAPB3_0_APBmslave0_PADDR[6], CoreAPB3_0_APBmslave0_PADDR[5], 
        CoreAPB3_0_APBmslave0_PADDR[4], CoreAPB3_0_APBmslave0_PADDR[3], 
        CoreAPB3_0_APBmslave0_PADDR[2], CoreAPB3_0_APBmslave0_PADDR[1], 
        CoreAPB3_0_APBmslave0_PADDR[0]}), .F_HM0_ENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .F_HM0_SEL(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc59, 
        nc60}), .F_HM0_TRANS1(), .F_HM0_WDATA({nc61, nc62, nc63, nc64, 
        nc65, nc66, nc67, nc68, nc69, nc70, nc71, nc72, nc73, nc74, 
        nc75, nc76, CoreAPB3_0_APBmslave0_PWDATA[15], 
        CoreAPB3_0_APBmslave0_PWDATA[14], 
        CoreAPB3_0_APBmslave0_PWDATA[13], 
        CoreAPB3_0_APBmslave0_PWDATA[12], 
        CoreAPB3_0_APBmslave0_PWDATA[11], 
        CoreAPB3_0_APBmslave0_PWDATA[10], 
        CoreAPB3_0_APBmslave0_PWDATA[9], 
        CoreAPB3_0_APBmslave0_PWDATA[8], 
        CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc77, nc78}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc79, nc80, nc81, nc82}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc83, nc84}), .FAB_XDATAOUT({nc85, nc86, nc87, nc88, nc89, 
        nc90, nc91, nc92}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc93, 
        nc94}), .FIC32_1_MASTER({nc95, nc96}), .FPGA_RESET_N(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), .H2F_INTERRUPT({
        nc97, nc98, nc99, nc100, nc101, nc102, nc103, nc104, nc105, 
        nc106, nc107, nc108, nc109, nc110, nc111, nc112}), .H2F_NMI(), 
        .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc113, nc114, nc115, nc116, nc117, nc118, 
        nc119, nc120, nc121, nc122, nc123, nc124, nc125, nc126}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc127, nc128, nc129, nc130, nc131, nc132, 
        nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, nc141, 
        nc142, nc143, nc144, nc145, nc146, nc147, nc148, nc149, nc150, 
        nc151, nc152, nc153, nc154, nc155, nc156, nc157, nc158}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc159, nc160, nc161, nc162, 
        nc163, nc164, nc165, nc166, nc167, nc168}), .TRACECLK(), 
        .TRACEDATA({nc169, nc170, nc171, nc172}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc173, nc174, nc175, 
        nc176}), .TXDF({nc177, nc178, nc179, nc180, nc181, nc182, 
        nc183, nc184}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc185, nc186, nc187, nc188})
        , .F_BRESP_HRESP0({nc189, nc190}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc191, nc192, nc193, nc194, nc195, nc196, 
        nc197, nc198, nc199, nc200, nc201, nc202, nc203, nc204, nc205, 
        nc206, nc207, nc208, nc209, nc210, nc211, nc212, nc213, nc214, 
        nc215, nc216, nc217, nc218, nc219, nc220, nc221, nc222, nc223, 
        nc224, nc225, nc226, nc227, nc228, nc229, nc230, nc231, nc232, 
        nc233, nc234, nc235, nc236, nc237, nc238, nc239, nc240, nc241, 
        nc242, nc243, nc244, nc245, nc246, nc247, nc248, nc249, nc250, 
        nc251, nc252, nc253, nc254}), .F_RID({nc255, nc256, nc257, 
        nc258}), .F_RLAST(), .F_RRESP_HRESP1({nc259, nc260}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc261, nc262, 
        nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, nc271, 
        nc272, nc273, nc274, nc275, nc276}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        CoreUARTapb_2_1_intr_or_2_Y, CoreUARTapb_2_0_intr_or_2_Y, 
        COREI2C_0_0_INT[0]}), .F2HCALIB(VCC_net_1), .F_DMAREADY({
        VCC_net_1, VCC_net_1}), .F_FM0_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(GND_net_1), 
        .F_FM0_READY(VCC_net_1), .F_FM0_SEL(GND_net_1), .F_FM0_SIZE({
        GND_net_1, GND_net_1}), .F_FM0_TRANS1(GND_net_1), .F_FM0_WDATA({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_FM0_WRITE(GND_net_1), .F_HM0_RDATA({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]}), .F_HM0_READY(
        VCC_net_1), .F_HM0_RESP(GND_net_1), .FAB_AVALID(VCC_net_1), 
        .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(LOCK), .FAB_RXACTIVE(VCC_net_1), 
        .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(GND_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(VCC_net_1), .XCLK_FAB(VCC_net_1), 
        .CLK_BASE(GL0_INST), .CLK_MDDR_APB(VCC_net_1), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), .SPI1_SCK_IN(
        GND_net_1), .SPI1_SDI_MGPIO11A_IN(GND_net_1), 
        .SPI1_SDO_MGPIO12A_IN(GND_net_1), .SPI1_SS0_MGPIO13A_IN(
        GND_net_1), .SPI1_SS1_MGPIO14A_IN(GND_net_1), 
        .SPI1_SS2_MGPIO15A_IN(GND_net_1), .SPI1_SS3_MGPIO16A_IN(
        GND_net_1), .SPI1_SS4_MGPIO17A_IN(GND_net_1), 
        .SPI1_SS5_MGPIO18A_IN(GND_net_1), .SPI1_SS6_MGPIO23A_IN(
        GND_net_1), .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc277, nc278, 
        nc279, nc280, nc281, nc282, nc283, nc284, nc285, nc286, nc287, 
        nc288, nc289, nc290, nc291, nc292}), .DRAM_BA({nc293, nc294, 
        nc295}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc296, nc297, nc298}), .DRAM_DQ_OUT({nc299, 
        nc300, nc301, nc302, nc303, nc304, nc305, nc306, nc307, nc308, 
        nc309, nc310, nc311, nc312, nc313, nc314, nc315, nc316}), 
        .DRAM_DQS_OUT({nc317, nc318, nc319}), .DRAM_FIFO_WE_OUT({nc320, 
        nc321}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc322, nc323, 
        nc324}), .DRAM_DQ_OE({nc325, nc326, nc327, nc328, nc329, nc330, 
        nc331, nc332, nc333, nc334, nc335, nc336, nc337, nc338, nc339, 
        nc340, nc341, nc342}), .DRAM_DQS_OE({nc343, nc344, nc345}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CCC_0_FCCC(
       GL0_INST,
       LOCK,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output GL0_INST;
output LOCK;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST_inst_1 (.A(GL0_net), .Y(GL0_INST));
    CCC #( .INIT(210'h0000007FB8000045164000318C6318C1F18C61EC0404040400101)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(LOCK), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module mss_sb_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb(
       TRIG_c,
       ECHO_c,
       PWM_c,
       COREI2C_0_0_SDA_IO,
       COREI2C_0_0_SCL_IO,
       DEVRST_N,
       BT_RX_c,
       BT_TX_c,
       GPS_RX_c,
       GPS_TX_c
    );
output [0:0] TRIG_c;
input  [1:1] ECHO_c;
output [10:1] PWM_c;
inout  COREI2C_0_0_SDA_IO;
inout  COREI2C_0_0_SCL_IO;
input  DEVRST_N;
output BT_RX_c;
input  BT_TX_c;
output GPS_RX_c;
input  GPS_TX_c;

    wire BIBUF_COREI2C_0_0_SDA_IO_Y, GND_net_1, 
        \COREI2C_0_0_SDAO_i[0] , BIBUF_COREI2C_0_0_SCL_IO_Y, 
        \COREI2C_0_0_SCLO_i[0] , SYSRESET_POR_net_1, 
        CoreUARTapb_2_1_intr_or_2_Y, CoreUARTapb_2_1_intr_or_1_Y, 
        CoreUARTapb_2_1_intr_or_0_Y, CoreUARTapb_2_1_RXRDY, 
        CoreUARTapb_2_1_TXRDY, CoreUARTapb_2_1_FRAMING_ERR, 
        CoreUARTapb_2_1_OVERFLOW, CoreUARTapb_2_1_PARITY_ERR, 
        CoreUARTapb_2_0_intr_or_2_Y, CoreUARTapb_2_0_intr_or_1_Y, 
        CoreUARTapb_2_0_intr_or_0_Y, CoreUARTapb_2_0_RXRDY, 
        CoreUARTapb_2_0_TXRDY, CoreUARTapb_2_0_FRAMING_ERR, 
        CoreUARTapb_2_0_OVERFLOW, CoreUARTapb_2_0_PARITY_ERR, GL0_INST, 
        LOCK, FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \iPSELS_0[4] , \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] , \iPSELS_0_0[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , \sercon[0] , \sercon[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , \serdat[0] , \serdat[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m_0[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m_1[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m_2[7] , 
        \CoreAPB3_0_APBmslave1_PRDATA_m[0] , 
        \CoreAPB3_0_APBmslave1_PRDATA_m[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] , 
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave3_PSELx, CoreAPB3_0_APBmslave2_PSELx, 
        CoreAPB3_0_APBmslave1_PSELx, CoreAPB3_0_APBmslave0_PSELx, 
        un4_PRDATA_1, controlReg14_3, r_N_4_mux, un12_PSELi, 
        un4_PRDATA, un1_PRDATA, PRDATA_regif_sn_N_39_mux, un14_PRDATA, 
        PRDATA_regif_sn_N_26, N_809, N_829, N_810, N_830, N_807, N_827, 
        N_808, N_828, N_812, N_832, N_806, N_826, N_813, N_833, N_811, 
        N_831, N_840, N_842, N_837, N_841, N_839, N_838, 
        \GPOUT_reg[1] , \CoreAPB3_0_APBmslave0_PWDATA[0] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , \gpin3_m_2_0[1] , 
        \gpin3_m[1] , MSS_HPMS_READY_int_RNI5CTC, GPOUT_reg40_2, 
        GPOUT_reg40, un1_WEn_1, \COREI2C_0_0_INT[0] , 
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , N_97_1, 
        CoreAPB3_0_APBmslave0_PENABLE, CoreAPB3_0_APBmslave0_PWRITE, 
        un1_WEn_0, \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[15] , un1_OEn_2, 
        un3_PRDATA_regif_1, psh_negedge_reg_1_sqmuxa_3_2, 
        controlReg24_3, mss_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, un1_OEn_1, 
        controlReg24_0, controlReg14_0, VCC_net_1;
    
    CoreAPB3_Z1 CoreAPB3_0 (.iPSELS_0({\iPSELS_0[4] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] }), .iPSELS_0_0({
        \iPSELS_0_0[4] }), .CoreAPB3_0_APBmslave2_PRDATA({
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_0({
        \CoreAPB3_0_APBmslave0_PRDATA_m_0[7] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_1({
        \CoreAPB3_0_APBmslave0_PRDATA_m_1[7] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2({
        \CoreAPB3_0_APBmslave0_PRDATA_m_2[7] }), 
        .CoreAPB3_0_APBmslave1_PRDATA_m({
        \CoreAPB3_0_APBmslave1_PRDATA_m[1] , 
        \CoreAPB3_0_APBmslave1_PRDATA_m[0] }), 
        .CoreAPB3_0_APBmslave4_PRDATA({
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] }), .sercon_0(
        \sercon[0] ), .sercon_2(\sercon[2] ), 
        .CoreAPB3_0_APBmslave0_PADDR_0(
        \CoreAPB3_0_APBmslave0_PADDR[0] ), 
        .CoreAPB3_0_APBmslave0_PADDR_7(
        \CoreAPB3_0_APBmslave0_PADDR[7] ), .serdat_0(\serdat[0] ), 
        .serdat_2(\serdat[2] ), .CoreAPB3_0_APBmslave0_PRDATA_m_0_d0(
        \CoreAPB3_0_APBmslave0_PRDATA_m[1] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_4(
        \CoreAPB3_0_APBmslave0_PRDATA_m[5] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_5(
        \CoreAPB3_0_APBmslave0_PRDATA_m[6] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_3(
        \CoreAPB3_0_APBmslave0_PRDATA_m[4] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2_d0(
        \CoreAPB3_0_APBmslave0_PRDATA_m[3] ), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_0_APBmslave2_PSELx(CoreAPB3_0_APBmslave2_PSELx), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .CoreAPB3_0_APBmslave0_PSELx(CoreAPB3_0_APBmslave0_PSELx), 
        .un4_PRDATA_1(un4_PRDATA_1), .controlReg14_3(controlReg14_3), 
        .r_N_4_mux(r_N_4_mux), .un12_PSELi(un12_PSELi), .un4_PRDATA(
        un4_PRDATA), .un1_PRDATA(un1_PRDATA), 
        .PRDATA_regif_sn_N_39_mux(PRDATA_regif_sn_N_39_mux), 
        .un14_PRDATA(un14_PRDATA), .PRDATA_regif_sn_N_26(
        PRDATA_regif_sn_N_26), .N_809(N_809), .N_829(N_829), .N_810(
        N_810), .N_830(N_830), .N_807(N_807), .N_827(N_827), .N_808(
        N_808), .N_828(N_828), .N_812(N_812), .N_832(N_832), .N_806(
        N_806), .N_826(N_826), .N_813(N_813), .N_833(N_833), .N_811(
        N_811), .N_831(N_831), .N_840(N_840), .N_842(N_842), .N_837(
        N_837), .N_841(N_841), .N_839(N_839), .N_838(N_838));
    BIBUF BIBUF_COREI2C_0_0_SDA_IO (.PAD(COREI2C_0_0_SDA_IO), .D(
        GND_net_1), .E(\COREI2C_0_0_SDAO_i[0] ), .Y(
        BIBUF_COREI2C_0_0_SDA_IO_Y));
    CoreGPIO_Z2 CoreGPIO_0_0 (.GPOUT_reg({\GPOUT_reg[1] }), .TRIG_c({
        TRIG_c[0]}), .CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .ECHO_c({ECHO_c[1]}), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] }), .gpin3_m_2_0({
        \gpin3_m_2_0[1] }), .gpin3_m({\gpin3_m[1] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .GPOUT_reg40_2(GPOUT_reg40_2), 
        .GPOUT_reg40(GPOUT_reg40), .un1_WEn_1(un1_WEn_1), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx));
    GND GND (.Y(GND_net_1));
    OR3 CoreUARTapb_2_1_intr_or_0 (.A(CoreUARTapb_2_1_FRAMING_ERR), .B(
        CoreUARTapb_2_1_OVERFLOW), .C(CoreUARTapb_2_1_PARITY_ERR), .Y(
        CoreUARTapb_2_1_intr_or_0_Y));
    OR3 CoreUARTapb_2_0_intr_or_1 (.A(CoreUARTapb_2_0_RXRDY), .B(
        CoreUARTapb_2_0_TXRDY), .C(GND_net_1), .Y(
        CoreUARTapb_2_0_intr_or_1_Y));
    COREI2C_Z3 COREI2C_0_0 (.COREI2C_0_0_SDAO_i({
        \COREI2C_0_0_SDAO_i[0] }), .COREI2C_0_0_SCLO_i({
        \COREI2C_0_0_SCLO_i[0] }), .COREI2C_0_0_INT({
        \COREI2C_0_0_INT[0] }), .CoreAPB3_0_APBmslave0_PADDR({
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_1({
        \CoreAPB3_0_APBmslave0_PRDATA_m_1[7] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_0({
        \CoreAPB3_0_APBmslave0_PRDATA_m_0[7] }), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2({
        \CoreAPB3_0_APBmslave0_PRDATA_m_2[7] }), .TRIG_c({TRIG_c[0]}), 
        .gpin3_m_2_0({\gpin3_m_2_0[1] }), .GPOUT_reg({\GPOUT_reg[1] }), 
        .gpin3_m({\gpin3_m[1] }), .CoreAPB3_0_APBmslave1_PRDATA_m({
        \CoreAPB3_0_APBmslave1_PRDATA_m[1] , 
        \CoreAPB3_0_APBmslave1_PRDATA_m[0] }), 
        .CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .sercon_0(\sercon[0] ), 
        .sercon_2(\sercon[2] ), .serdat_2(\serdat[2] ), .serdat_0(
        \serdat[0] ), .CoreAPB3_0_APBmslave0_PRDATA_m_0_d0(
        \CoreAPB3_0_APBmslave0_PRDATA_m[1] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_4(
        \CoreAPB3_0_APBmslave0_PRDATA_m[5] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_2_d0(
        \CoreAPB3_0_APBmslave0_PRDATA_m[3] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_3(
        \CoreAPB3_0_APBmslave0_PRDATA_m[4] ), 
        .CoreAPB3_0_APBmslave0_PRDATA_m_5(
        \CoreAPB3_0_APBmslave0_PRDATA_m[6] ), .un12_PSELi(un12_PSELi), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .r_N_4_mux(r_N_4_mux), .N_97_1(N_97_1), 
        .controlReg14_3(controlReg14_3), .un4_PRDATA_1(un4_PRDATA_1), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .un1_WEn_1(un1_WEn_1), .BIBUF_COREI2C_0_0_SCL_IO_Y(
        BIBUF_COREI2C_0_0_SCL_IO_Y), .BIBUF_COREI2C_0_0_SDA_IO_Y(
        BIBUF_COREI2C_0_0_SDA_IO_Y), .un1_WEn_0(un1_WEn_0), 
        .un14_PRDATA(un14_PRDATA), .un1_PRDATA(un1_PRDATA), 
        .un4_PRDATA(un4_PRDATA), .CoreAPB3_0_APBmslave0_PSELx(
        CoreAPB3_0_APBmslave0_PSELx), .GPOUT_reg40_2(GPOUT_reg40_2), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .GPOUT_reg40(GPOUT_reg40));
    CoreResetP_Z7 CORERESETP_0 (.MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .SYSRESET_POR(SYSRESET_POR_net_1), 
        .mss_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), 
        .mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    OR3 CoreUARTapb_2_0_intr_or_2 (.A(CoreUARTapb_2_0_intr_or_1_Y), .B(
        CoreUARTapb_2_0_intr_or_0_Y), .C(GND_net_1), .Y(
        CoreUARTapb_2_0_intr_or_2_Y));
    OR3 CoreUARTapb_2_0_intr_or_0 (.A(CoreUARTapb_2_0_FRAMING_ERR), .B(
        CoreUARTapb_2_0_OVERFLOW), .C(CoreUARTapb_2_0_PARITY_ERR), .Y(
        CoreUARTapb_2_0_intr_or_0_Y));
    mss_sb_CoreUARTapb_2_0_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s 
        CoreUARTapb_2_0 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PRDATA({
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .un1_OEn_2(un1_OEn_2), .controlReg24_3(
        controlReg24_3), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .un1_OEn_1(un1_OEn_1), 
        .controlReg24_0(controlReg24_0), .controlReg14_3(
        controlReg14_3), .controlReg14_0(controlReg14_0), 
        .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR), 
        .N_97_1(N_97_1), .CoreAPB3_0_APBmslave2_PSELx(
        CoreAPB3_0_APBmslave2_PSELx), .psh_negedge_reg_1_sqmuxa_3_2(
        psh_negedge_reg_1_sqmuxa_3_2), .CoreUARTapb_2_0_FRAMING_ERR(
        CoreUARTapb_2_0_FRAMING_ERR), .CoreUARTapb_2_0_OVERFLOW(
        CoreUARTapb_2_0_OVERFLOW), .CoreUARTapb_2_0_RXRDY(
        CoreUARTapb_2_0_RXRDY), .CoreUARTapb_2_0_TXRDY(
        CoreUARTapb_2_0_TXRDY), .un1_WEn_1(un1_WEn_1), .un1_WEn_0(
        un1_WEn_0), .BT_RX_c(BT_RX_c), .BT_TX_c(BT_TX_c));
    mss_sb_CoreUARTapb_2_1_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s 
        CoreUARTapb_2_1 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .un3_PRDATA_regif_1(un3_PRDATA_regif_1), 
        .CoreUARTapb_2_1_PARITY_ERR(CoreUARTapb_2_1_PARITY_ERR), 
        .N_97_1(N_97_1), .CoreUARTapb_2_1_RXRDY(CoreUARTapb_2_1_RXRDY), 
        .CoreUARTapb_2_1_TXRDY(CoreUARTapb_2_1_TXRDY), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .controlReg14_0(controlReg14_0), .controlReg24_0(
        controlReg24_0), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .psh_negedge_reg_1_sqmuxa_3_2(
        psh_negedge_reg_1_sqmuxa_3_2), .CoreUARTapb_2_1_FRAMING_ERR(
        CoreUARTapb_2_1_FRAMING_ERR), .CoreUARTapb_2_1_OVERFLOW(
        CoreUARTapb_2_1_OVERFLOW), .un1_WEn_1(un1_WEn_1), .un1_WEn_0(
        un1_WEn_0), .un1_OEn_2(un1_OEn_2), .un1_OEn_1(un1_OEn_1), 
        .GPS_RX_c(GPS_RX_c), .GPS_TX_c(GPS_TX_c));
    OR3 CoreUARTapb_2_1_intr_or_2 (.A(CoreUARTapb_2_1_intr_or_1_Y), .B(
        CoreUARTapb_2_1_intr_or_0_Y), .C(GND_net_1), .Y(
        CoreUARTapb_2_1_intr_or_2_Y));
    corepwm_Z5 corepwm_0_0 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .iPSELS_0_0({
        \iPSELS_0_0[4] }), .iPSELS_0({\iPSELS_0[4] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .CoreAPB3_0_APBmslave4_PRDATA({
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] }), .PWM_c({PWM_c[10], 
        PWM_c[9], PWM_c[8], PWM_c[7], PWM_c[6], PWM_c[5], PWM_c[4], 
        PWM_c[3], PWM_c[2], PWM_c[1]}), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .N_97_1(N_97_1), .controlReg14_3(controlReg14_3), 
        .PRDATA_regif_sn_N_26(PRDATA_regif_sn_N_26), .N_842(N_842), 
        .N_841(N_841), .N_840(N_840), .un1_OEn_2(un1_OEn_2), 
        .un3_PRDATA_regif_1(un3_PRDATA_regif_1), 
        .psh_negedge_reg_1_sqmuxa_3_2(psh_negedge_reg_1_sqmuxa_3_2), 
        .N_813(N_813), .N_811(N_811), .N_806(N_806), .N_812(N_812), 
        .N_807(N_807), .N_808(N_808), .N_810(N_810), .N_809(N_809), 
        .controlReg24_3(controlReg24_3), .PRDATA_regif_sn_N_39_mux(
        PRDATA_regif_sn_N_39_mux), .N_833(N_833), .N_831(N_831), 
        .N_828(N_828), .N_826(N_826), .N_832(N_832), .N_827(N_827), 
        .N_830(N_830), .N_829(N_829), .N_837(N_837), .N_839(N_839), 
        .N_838(N_838));
    mss_sb_MSS mss_sb_MSS_0 (.CoreAPB3_0_APBmslave0_PADDR({
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] }), 
        .CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .COREI2C_0_0_INT({
        \COREI2C_0_0_INT[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .mss_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), 
        .CoreUARTapb_2_0_intr_or_2_Y(CoreUARTapb_2_0_intr_or_2_Y), 
        .CoreUARTapb_2_1_intr_or_2_Y(CoreUARTapb_2_1_intr_or_2_Y), 
        .LOCK(LOCK), .GL0_INST(GL0_INST));
    VCC VCC (.Y(VCC_net_1));
    mss_sb_CCC_0_FCCC CCC_0 (.GL0_INST(GL0_INST), .LOCK(LOCK), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    BIBUF BIBUF_COREI2C_0_0_SCL_IO (.PAD(COREI2C_0_0_SCL_IO), .D(
        GND_net_1), .E(\COREI2C_0_0_SCLO_i[0] ), .Y(
        BIBUF_COREI2C_0_0_SCL_IO_Y));
    mss_sb_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    OR3 CoreUARTapb_2_1_intr_or_1 (.A(CoreUARTapb_2_1_RXRDY), .B(
        CoreUARTapb_2_1_TXRDY), .C(GND_net_1), .Y(
        CoreUARTapb_2_1_intr_or_1_Y));
    
endmodule


module mss(
       ECHO,
       PWM,
       TRIG,
       BT_TX,
       DEVRST_N,
       GPS_TX,
       BT_RX,
       GPS_RX,
       COREI2C_0_0_SCL_IO,
       COREI2C_0_0_SDA_IO
    );
input  [1:0] ECHO;
output [10:1] PWM;
output [1:0] TRIG;
input  BT_TX;
input  DEVRST_N;
input  GPS_TX;
output BT_RX;
output GPS_RX;
inout  COREI2C_0_0_SCL_IO;
inout  COREI2C_0_0_SDA_IO;

    wire VCC_net_1, GND_net_1, BT_TX_c, \ECHO_c[1] , GPS_TX_c, BT_RX_c, 
        GPS_RX_c, \PWM_c[1] , \PWM_c[2] , \PWM_c[3] , \PWM_c[4] , 
        \PWM_c[5] , \PWM_c[6] , \PWM_c[7] , \PWM_c[8] , \PWM_c[9] , 
        \PWM_c[10] , \TRIG_c[0] ;
    
    OUTBUF BT_RX_obuf (.D(BT_RX_c), .PAD(BT_RX));
    OUTBUF \PWM_obuf[3]  (.D(\PWM_c[3] ), .PAD(PWM[3]));
    mss_sb mss_sb_0 (.TRIG_c({\TRIG_c[0] }), .ECHO_c({\ECHO_c[1] }), 
        .PWM_c({\PWM_c[10] , \PWM_c[9] , \PWM_c[8] , \PWM_c[7] , 
        \PWM_c[6] , \PWM_c[5] , \PWM_c[4] , \PWM_c[3] , \PWM_c[2] , 
        \PWM_c[1] }), .COREI2C_0_0_SDA_IO(COREI2C_0_0_SDA_IO), 
        .COREI2C_0_0_SCL_IO(COREI2C_0_0_SCL_IO), .DEVRST_N(DEVRST_N), 
        .BT_RX_c(BT_RX_c), .BT_TX_c(BT_TX_c), .GPS_RX_c(GPS_RX_c), 
        .GPS_TX_c(GPS_TX_c));
    GND GND (.Y(GND_net_1));
    INBUF \ECHO_ibuf[1]  (.PAD(ECHO[1]), .Y(\ECHO_c[1] ));
    OUTBUF \PWM_obuf[7]  (.D(\PWM_c[7] ), .PAD(PWM[7]));
    OUTBUF GPS_RX_obuf (.D(GPS_RX_c), .PAD(GPS_RX));
    OUTBUF \TRIG_obuf[0]  (.D(\TRIG_c[0] ), .PAD(TRIG[0]));
    OUTBUF \PWM_obuf[1]  (.D(\PWM_c[1] ), .PAD(PWM[1]));
    OUTBUF \PWM_obuf[10]  (.D(\PWM_c[10] ), .PAD(PWM[10]));
    OUTBUF \PWM_obuf[2]  (.D(\PWM_c[2] ), .PAD(PWM[2]));
    INBUF BT_TX_ibuf (.PAD(BT_TX), .Y(BT_TX_c));
    OUTBUF \PWM_obuf[9]  (.D(\PWM_c[9] ), .PAD(PWM[9]));
    OUTBUF \PWM_obuf[6]  (.D(\PWM_c[6] ), .PAD(PWM[6]));
    OUTBUF \PWM_obuf[8]  (.D(\PWM_c[8] ), .PAD(PWM[8]));
    INBUF GPS_TX_ibuf (.PAD(GPS_TX), .Y(GPS_TX_c));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF \PWM_obuf[4]  (.D(\PWM_c[4] ), .PAD(PWM[4]));
    OUTBUF \TRIG_obuf[1]  (.D(GND_net_1), .PAD(TRIG[1]));
    OUTBUF \PWM_obuf[5]  (.D(\PWM_c[5] ), .PAD(PWM[5]));
    
endmodule
