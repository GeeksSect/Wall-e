`timescale 1 ns/100 ps
// Version: v11.6 SP1 11.6.1.6


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module RCOSC_1MHZ(
       CLKOUT
    );
output CLKOUT;

    
endmodule


module COREAPB3_MUXPTOB3(
       period_reg,
       pwm_enable_reg,
       PRDATA_regif_0_0,
       sersta_m_0,
       PRDATA_regif_9_i_0,
       PRDATA_regif_9_i_1,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR,
       CoreAPB3_0_APBmslave4_PRDATA,
       PRDATA_regif_12_0,
       sersta_m,
       serdat_m,
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave2_PRDATA,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR_3,
       CoreAPB3_0_APBmslave0_PADDR_2,
       CoreAPB3_0_APBmslave0_PADDR_0,
       CoreAPB3_0_APBmslave0_PADDR_5,
       serdat_4,
       serdat_0,
       \PRDATAi[0]_2 ,
       \PRDATAi[0]_0 ,
       \PRDATAi[0]_6 ,
       \PRDATAi[0]_1 ,
       \PRDATAi[0]_4 ,
       sercon_m_4,
       sercon_m_0,
       sercon_m_6,
       CoreAPB3_0_APBmslave4_PSELx,
       N_513,
       N_699,
       N_428,
       N_529,
       N_411,
       un12_PSELi,
       un9_PRDATA_2_0,
       psh_enable_reg1_1_sqmuxa_0,
       N_629,
       CoreAPB3_0_APBmslave1_PSELx,
       CoreAPB3_0_APBmslave3_PSELx,
       N_426,
       N_432,
       N_685,
       N_680,
       N_684,
       N_681,
       N_703,
       N_698,
       N_702,
       N_691,
       CoreAPB3_0_APBmslave0_PSELx,
       N_709,
       N_679,
       N_678,
       N_506,
       N_711,
       N_140,
       N_710,
       un4_PRDATA,
       N_700,
       N_687,
       N_705,
       N_688,
       N_706,
       N_690,
       N_708,
       N_689,
       N_707,
       N_686,
       N_704,
       PRDATA_regif_sn_N_20_i_1,
       N_660
    );
input  [5:5] period_reg;
input  [6:6] pwm_enable_reg;
input  [5:5] PRDATA_regif_0_0;
input  [1:1] sersta_m_0;
input  [4:4] PRDATA_regif_9_i_0;
input  [4:4] PRDATA_regif_9_i_1;
input  [14:12] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR;
input  [7:0] CoreAPB3_0_APBmslave4_PRDATA;
input  [1:1] PRDATA_regif_12_0;
input  [3:3] sersta_m;
input  [6:6] serdat_m;
input  [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave2_PRDATA;
output [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
input  CoreAPB3_0_APBmslave0_PADDR_3;
input  CoreAPB3_0_APBmslave0_PADDR_2;
input  CoreAPB3_0_APBmslave0_PADDR_0;
input  CoreAPB3_0_APBmslave0_PADDR_5;
input  serdat_4;
input  serdat_0;
input  \PRDATAi[0]_2 ;
input  \PRDATAi[0]_0 ;
input  \PRDATAi[0]_6 ;
input  \PRDATAi[0]_1 ;
input  \PRDATAi[0]_4 ;
input  sercon_m_4;
input  sercon_m_0;
input  sercon_m_6;
input  CoreAPB3_0_APBmslave4_PSELx;
input  N_513;
input  N_699;
input  N_428;
input  N_529;
input  N_411;
input  un12_PSELi;
input  un9_PRDATA_2_0;
input  psh_enable_reg1_1_sqmuxa_0;
input  N_629;
input  CoreAPB3_0_APBmslave1_PSELx;
input  CoreAPB3_0_APBmslave3_PSELx;
input  N_426;
output N_432;
input  N_685;
input  N_680;
input  N_684;
input  N_681;
input  N_703;
input  N_698;
input  N_702;
input  N_691;
input  CoreAPB3_0_APBmslave0_PSELx;
input  N_709;
input  N_679;
input  N_678;
input  N_506;
input  N_711;
input  N_140;
input  N_710;
input  un4_PRDATA;
input  N_700;
input  N_687;
input  N_705;
input  N_688;
input  N_706;
input  N_690;
input  N_708;
input  N_689;
input  N_707;
input  N_686;
input  N_704;
input  PRDATA_regif_sn_N_20_i_1;
input  N_660;

    wire \PRDATA_5_d[3]_net_1 , N_108, \PRDATA_5_1_1[5]_net_1 , 
        \PRDATA_5_1[5]_net_1 , N_110, \PRDATA_4_bm_1[4]_net_1 , 
        \PRDATA_4_bm[4]_net_1 , \PRDATA_5_d_1[4]_net_1 , 
        \PRDATA_5_d[4]_net_1 , \PRDATA_4_s[3]_net_1 , 
        \PRDATA_4_ns_1[3]_net_1 , N_100, \PRDATA_4_am[4]_net_1 , N_101, 
        \PRDATA_4_am[6]_net_1 , \PRDATA_4_bm[6]_net_1 , N_103, 
        \PRDATA_4_am[0]_net_1 , \PRDATA_4_bm[0]_net_1 , N_97, 
        \PRDATA_5_s[3]_net_1 , \PRDATA_5_d[7]_net_1 , 
        \PRDATA_5_d[2]_net_1 , \PRDATA_5_d[6]_net_1 , PRDATA_sn_N_5, 
        \PRDATA_4_d[1]_net_1 , \PRDATA_4_d[7]_net_1 , 
        \PRDATA_4_d[2]_net_1 , \PRDATA_4_d[5]_net_1 , N_112, N_107, 
        N_111, \PRDATA_5_d[1]_net_1 , \PRDATA_5_d[0]_net_1 , 
        PRDATA_sn_N_9_mux, N_98, N_109, N_106, N_105, N_104, N_99, 
        N_102, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h0D0F) )  \PRDATA_5_1[5]  (.A(N_428), .B(N_529), 
        .C(N_411), .D(\PRDATA_5_1_1[5]_net_1 ), .Y(
        \PRDATA_5_1[5]_net_1 ));
    CFG4 #( .INIT(16'hF0DD) )  \PRDATA_5[5]  (.A(\PRDATA_5_1[5]_net_1 )
        , .B(PRDATA_regif_0_0[5]), .C(CoreAPB3_0_APBmslave4_PRDATA[5]), 
        .D(CoreAPB3_0_APBmslave4_PSELx), .Y(N_110));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[1]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[1]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_679), .Y(
        \PRDATA_5_d[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \PRDATA_4_ns[0]  (.A(\PRDATA_4_s[3]_net_1 )
        , .B(\PRDATA_4_am[0]_net_1 ), .C(\PRDATA_4_bm[0]_net_1 ), .Y(
        N_97));
    CFG2 #( .INIT(4'h2) )  \PRDATA_5_s[3]  (.A(N_513), .B(
        CoreAPB3_0_APBmslave4_PSELx), .Y(\PRDATA_5_s[3]_net_1 ));
    CFG4 #( .INIT(16'h0AC0) )  \PRDATA_5_1_1[5]  (.A(period_reg[5]), 
        .B(pwm_enable_reg[6]), .C(CoreAPB3_0_APBmslave0_PADDR_3), .D(
        CoreAPB3_0_APBmslave0_PADDR_2), .Y(\PRDATA_5_1_1[5]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[6]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[6]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_684), .Y(
        \PRDATA_5_d[6]_net_1 ));
    CFG4 #( .INIT(16'hB010) )  \PRDATA[14]  (.A(N_513), .B(N_140), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_710), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14]));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_am[0]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[0]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[0]), .Y(\PRDATA_4_am[0]_net_1 ));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[4]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_109), .D(N_101), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4]));
    CFG3 #( .INIT(8'hE4) )  \PRDATA_5[7]  (.A(\PRDATA_5_s[3]_net_1 ), 
        .B(\PRDATA_5_d[7]_net_1 ), .C(N_703), .Y(N_112));
    CFG4 #( .INIT(16'hAA02) )  \PRDATA_4_bm[4]  (.A(un12_PSELi), .B(
        CoreAPB3_0_APBmslave0_PADDR_0), .C(\PRDATA_4_bm_1[4]_net_1 ), 
        .D(sercon_m_4), .Y(\PRDATA_4_bm[4]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[10]  (.A(N_513), .B(N_688), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_706), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10]));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[2]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_107), .D(N_99), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_d[1]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[1]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[1]), .Y(\PRDATA_4_d[1]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[0]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[0]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_678), .Y(
        \PRDATA_5_d[0]_net_1 ));
    CFG4 #( .INIT(16'h0E1F) )  \PRDATA_4_ns_1[3]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[3]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[3]), .Y(\PRDATA_4_ns_1[3]_net_1 ));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[1]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_106), .D(N_98), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_4_ns[4]  (.A(
        \PRDATA_4_am[4]_net_1 ), .B(\PRDATA_4_s[3]_net_1 ), .C(
        \PRDATA_4_bm[4]_net_1 ), .Y(N_101));
    CFG4 #( .INIT(16'h1F5F) )  \PRDATA_4_bm_1[4]  (.A(sersta_m_0[1]), 
        .B(serdat_4), .C(un9_PRDATA_2_0), .D(
        psh_enable_reg1_1_sqmuxa_0), .Y(\PRDATA_4_bm_1[4]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[8]  (.A(N_513), .B(N_686), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_704), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8]));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_4_ns[6]  (.A(
        \PRDATA_4_am[6]_net_1 ), .B(\PRDATA_4_s[3]_net_1 ), .C(
        \PRDATA_4_bm[6]_net_1 ), .Y(N_103));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[12]  (.A(N_513), .B(N_690), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_708), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12]));
    CFG4 #( .INIT(16'h8F80) )  \PRDATA_5[1]  (.A(PRDATA_regif_12_0[1]), 
        .B(PRDATA_regif_sn_N_20_i_1), .C(\PRDATA_5_s[3]_net_1 ), .D(
        \PRDATA_5_d[1]_net_1 ), .Y(N_106));
    CFG3 #( .INIT(8'hE4) )  \PRDATA_5[2]  (.A(\PRDATA_5_s[3]_net_1 ), 
        .B(\PRDATA_5_d[2]_net_1 ), .C(N_698), .Y(N_107));
    CFG4 #( .INIT(16'hD580) )  \PRDATA_4[7]  (.A(\PRDATA_4_s[3]_net_1 )
        , .B(un12_PSELi), .C(\PRDATAi[0]_6 ), .D(\PRDATA_4_d[7]_net_1 )
        , .Y(N_104));
    CFG4 #( .INIT(16'hCCC8) )  \PRDATA_4_bm[6]  (.A(sersta_m[3]), .B(
        un12_PSELi), .C(serdat_m[6]), .D(sercon_m_6), .Y(
        \PRDATA_4_bm[6]_net_1 ));
    CFG4 #( .INIT(16'h3F2E) )  \PRDATA_5_d_1[4]  (.A(
        PRDATA_regif_9_i_0[4]), .B(CoreAPB3_0_APBmslave0_PADDR_5), .C(
        N_629), .D(PRDATA_regif_9_i_1[4]), .Y(\PRDATA_5_d_1[4]_net_1 ));
    CFG4 #( .INIT(16'hD580) )  \PRDATA_4[5]  (.A(\PRDATA_4_s[3]_net_1 )
        , .B(un12_PSELi), .C(\PRDATAi[0]_4 ), .D(\PRDATA_4_d[5]_net_1 )
        , .Y(N_102));
    CFG4 #( .INIT(16'h5140) )  \PRDATA[5]  (.A(PRDATA_sn_N_9_mux), .B(
        PRDATA_sn_N_5), .C(N_110), .D(N_102), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5]));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hB1) )  \PRDATA_5_d[4]  (.A(
        CoreAPB3_0_APBmslave4_PSELx), .B(\PRDATA_5_d_1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave4_PRDATA[4]), .Y(\PRDATA_5_d[4]_net_1 ));
    CFG4 #( .INIT(16'h8F80) )  \PRDATA_5[0]  (.A(N_660), .B(
        PRDATA_regif_sn_N_20_i_1), .C(\PRDATA_5_s[3]_net_1 ), .D(
        \PRDATA_5_d[0]_net_1 ), .Y(N_105));
    CFG4 #( .INIT(16'hD580) )  \PRDATA_4[1]  (.A(\PRDATA_4_s[3]_net_1 )
        , .B(un12_PSELi), .C(\PRDATAi[0]_0 ), .D(\PRDATA_4_d[1]_net_1 )
        , .Y(N_98));
    CFG4 #( .INIT(16'hB010) )  \PRDATA[15]  (.A(N_513), .B(N_506), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_711), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15]));
    CFG4 #( .INIT(16'hAFBF) )  PRDATA_sn_m4 (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(PRDATA_sn_N_5)
        );
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[7]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[7]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_685), .Y(
        \PRDATA_5_d[7]_net_1 ));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_am[4]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[4]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[4]), .Y(\PRDATA_4_am[4]_net_1 ));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[0]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_105), .D(N_97), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]));
    CFG4 #( .INIT(16'hF4B0) )  \PRDATA_5[3]  (.A(
        CoreAPB3_0_APBmslave4_PSELx), .B(N_513), .C(
        \PRDATA_5_d[3]_net_1 ), .D(N_699), .Y(N_108));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[3]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_108), .D(N_100), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3]));
    CFG4 #( .INIT(16'hAF8F) )  PRDATA_sn_m7 (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        PRDATA_sn_N_9_mux));
    CFG3 #( .INIT(8'hE4) )  \PRDATA_5[4]  (.A(\PRDATA_5_s[3]_net_1 ), 
        .B(\PRDATA_5_d[4]_net_1 ), .C(N_700), .Y(N_109));
    CFG4 #( .INIT(16'h0040) )  \PSELSBUS_0_a2[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(N_432));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_d[7]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[7]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[7]), .Y(\PRDATA_4_d[7]_net_1 ));
    CFG4 #( .INIT(16'h8B03) )  \PRDATA_4_ns[3]  (.A(un12_PSELi), .B(
        \PRDATA_4_s[3]_net_1 ), .C(\PRDATA_4_ns_1[3]_net_1 ), .D(
        \PRDATAi[0]_2 ), .Y(N_100));
    CFG4 #( .INIT(16'hC8C0) )  \PRDATA_4_bm[0]  (.A(serdat_0), .B(
        un12_PSELi), .C(sercon_m_0), .D(un4_PRDATA), .Y(
        \PRDATA_4_bm[0]_net_1 ));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_d[5]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[5]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[5]), .Y(\PRDATA_4_d[5]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[9]  (.A(N_513), .B(N_687), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_705), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9]));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[6]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_111), .D(N_103), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6]));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[13]  (.A(N_513), .B(N_691), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_709), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13]));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_am[6]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[6]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[6]), .Y(\PRDATA_4_am[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[2]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[2]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_680), .Y(
        \PRDATA_5_d[2]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_5_d[3]  (.A(
        CoreAPB3_0_APBmslave4_PRDATA[3]), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(N_681), .Y(
        \PRDATA_5_d[3]_net_1 ));
    CFG4 #( .INIT(16'hF1E0) )  \PRDATA_4_d[2]  (.A(
        CoreAPB3_0_APBmslave1_PSELx), .B(CoreAPB3_0_APBmslave3_PSELx), 
        .C(CoreAPB3_0_APBmslave3_PRDATA[2]), .D(
        CoreAPB3_0_APBmslave2_PRDATA[2]), .Y(\PRDATA_4_d[2]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \PRDATA_5[6]  (.A(\PRDATA_5_s[3]_net_1 ), 
        .B(\PRDATA_5_d[6]_net_1 ), .C(N_702), .Y(N_111));
    CFG4 #( .INIT(16'hD580) )  \PRDATA_4[2]  (.A(\PRDATA_4_s[3]_net_1 )
        , .B(un12_PSELi), .C(\PRDATAi[0]_1 ), .D(\PRDATA_4_d[2]_net_1 )
        , .Y(N_99));
    CFG4 #( .INIT(16'h3120) )  \PRDATA[7]  (.A(PRDATA_sn_N_5), .B(
        PRDATA_sn_N_9_mux), .C(N_112), .D(N_104), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7]));
    CFG4 #( .INIT(16'h1000) )  \PRDATA_4_s[3]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        \PRDATA_4_s[3]_net_1 ));
    CFG4 #( .INIT(16'hE040) )  \PRDATA[11]  (.A(N_513), .B(N_689), .C(
        CoreAPB3_0_APBmslave0_PSELx), .D(N_707), .Y(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11]));
    
endmodule


module CoreAPB3_Z1_layer0(
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR,
       period_reg,
       pwm_enable_reg,
       PRDATA_regif_0_0,
       sersta_m_0,
       PRDATA_regif_9_i_0,
       PRDATA_regif_9_i_1,
       CoreAPB3_0_APBmslave4_PRDATA,
       PRDATA_regif_12_0,
       sersta_m,
       serdat_m,
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave2_PRDATA,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR_3,
       CoreAPB3_0_APBmslave0_PADDR_2,
       CoreAPB3_0_APBmslave0_PADDR_0,
       CoreAPB3_0_APBmslave0_PADDR_5,
       serdat_4,
       serdat_0,
       \PRDATAi[0]_2 ,
       \PRDATAi[0]_0 ,
       \PRDATAi[0]_6 ,
       \PRDATAi[0]_1 ,
       \PRDATAi[0]_4 ,
       sercon_m_4,
       sercon_m_0,
       sercon_m_6,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave0_PSELx,
       CoreAPB3_0_APBmslave4_PSELx,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_0_APBmslave1_PSELx,
       N_513,
       N_699,
       N_428,
       N_529,
       N_411,
       un12_PSELi,
       un9_PRDATA_2_0,
       psh_enable_reg1_1_sqmuxa_0,
       N_629,
       N_432,
       N_685,
       N_680,
       N_684,
       N_681,
       N_703,
       N_698,
       N_702,
       N_691,
       N_709,
       N_679,
       N_678,
       N_506,
       N_711,
       N_140,
       N_710,
       un4_PRDATA,
       N_700,
       N_687,
       N_705,
       N_688,
       N_706,
       N_690,
       N_708,
       N_689,
       N_707,
       N_686,
       N_704,
       PRDATA_regif_sn_N_20_i_1,
       N_660
    );
input  [15:12] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR;
input  [5:5] period_reg;
input  [6:6] pwm_enable_reg;
input  [5:5] PRDATA_regif_0_0;
input  [1:1] sersta_m_0;
input  [4:4] PRDATA_regif_9_i_0;
input  [4:4] PRDATA_regif_9_i_1;
input  [7:0] CoreAPB3_0_APBmslave4_PRDATA;
input  [1:1] PRDATA_regif_12_0;
input  [3:3] sersta_m;
input  [6:6] serdat_m;
input  [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave2_PRDATA;
output [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
input  CoreAPB3_0_APBmslave0_PADDR_3;
input  CoreAPB3_0_APBmslave0_PADDR_2;
input  CoreAPB3_0_APBmslave0_PADDR_0;
input  CoreAPB3_0_APBmslave0_PADDR_5;
input  serdat_4;
input  serdat_0;
input  \PRDATAi[0]_2 ;
input  \PRDATAi[0]_0 ;
input  \PRDATAi[0]_6 ;
input  \PRDATAi[0]_1 ;
input  \PRDATAi[0]_4 ;
input  sercon_m_4;
input  sercon_m_0;
input  sercon_m_6;
input  mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave0_PSELx;
output CoreAPB3_0_APBmslave4_PSELx;
output CoreAPB3_0_APBmslave3_PSELx;
output CoreAPB3_0_APBmslave1_PSELx;
input  N_513;
input  N_699;
input  N_428;
input  N_529;
input  N_411;
input  un12_PSELi;
input  un9_PRDATA_2_0;
input  psh_enable_reg1_1_sqmuxa_0;
input  N_629;
output N_432;
input  N_685;
input  N_680;
input  N_684;
input  N_681;
input  N_703;
input  N_698;
input  N_702;
input  N_691;
input  N_709;
input  N_679;
input  N_678;
input  N_506;
input  N_711;
input  N_140;
input  N_710;
input  un4_PRDATA;
input  N_700;
input  N_687;
input  N_705;
input  N_688;
input  N_706;
input  N_690;
input  N_708;
input  N_689;
input  N_707;
input  N_686;
input  N_704;
input  PRDATA_regif_sn_N_20_i_1;
input  N_660;

    wire N_426, GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h4000) )  \iPSELS_0_a2[3]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave3_PSELx));
    CFG4 #( .INIT(16'h1000) )  \iPSELS[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave1_PSELx));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0020) )  \iPSELS_0_RNI7Q8I1[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave4_PSELx));
    COREAPB3_MUXPTOB3 u_mux_p_to_b3 (.period_reg({period_reg[5]}), 
        .pwm_enable_reg({pwm_enable_reg[6]}), .PRDATA_regif_0_0({
        PRDATA_regif_0_0[5]}), .sersta_m_0({sersta_m_0[1]}), 
        .PRDATA_regif_9_i_0({PRDATA_regif_9_i_0[4]}), 
        .PRDATA_regif_9_i_1({PRDATA_regif_9_i_1[4]}), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR({
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]}), 
        .CoreAPB3_0_APBmslave4_PRDATA({CoreAPB3_0_APBmslave4_PRDATA[7], 
        CoreAPB3_0_APBmslave4_PRDATA[6], 
        CoreAPB3_0_APBmslave4_PRDATA[5], 
        CoreAPB3_0_APBmslave4_PRDATA[4], 
        CoreAPB3_0_APBmslave4_PRDATA[3], 
        CoreAPB3_0_APBmslave4_PRDATA[2], 
        CoreAPB3_0_APBmslave4_PRDATA[1], 
        CoreAPB3_0_APBmslave4_PRDATA[0]}), .PRDATA_regif_12_0({
        PRDATA_regif_12_0[1]}), .sersta_m({sersta_m[3]}), .serdat_m({
        serdat_m[6]}), .CoreAPB3_0_APBmslave3_PRDATA({
        CoreAPB3_0_APBmslave3_PRDATA[7], 
        CoreAPB3_0_APBmslave3_PRDATA[6], 
        CoreAPB3_0_APBmslave3_PRDATA[5], 
        CoreAPB3_0_APBmslave3_PRDATA[4], 
        CoreAPB3_0_APBmslave3_PRDATA[3], 
        CoreAPB3_0_APBmslave3_PRDATA[2], 
        CoreAPB3_0_APBmslave3_PRDATA[1], 
        CoreAPB3_0_APBmslave3_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave2_PRDATA({CoreAPB3_0_APBmslave2_PRDATA[7], 
        CoreAPB3_0_APBmslave2_PRDATA[6], 
        CoreAPB3_0_APBmslave2_PRDATA[5], 
        CoreAPB3_0_APBmslave2_PRDATA[4], 
        CoreAPB3_0_APBmslave2_PRDATA[3], 
        CoreAPB3_0_APBmslave2_PRDATA[2], 
        CoreAPB3_0_APBmslave2_PRDATA[1], 
        CoreAPB3_0_APBmslave2_PRDATA[0]}), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave0_PADDR_3(CoreAPB3_0_APBmslave0_PADDR_3), 
        .CoreAPB3_0_APBmslave0_PADDR_2(CoreAPB3_0_APBmslave0_PADDR_2), 
        .CoreAPB3_0_APBmslave0_PADDR_0(CoreAPB3_0_APBmslave0_PADDR_0), 
        .CoreAPB3_0_APBmslave0_PADDR_5(CoreAPB3_0_APBmslave0_PADDR_5), 
        .serdat_4(serdat_4), .serdat_0(serdat_0), .\PRDATAi[0]_2 (
        \PRDATAi[0]_2 ), .\PRDATAi[0]_0 (\PRDATAi[0]_0 ), 
        .\PRDATAi[0]_6 (\PRDATAi[0]_6 ), .\PRDATAi[0]_1 (
        \PRDATAi[0]_1 ), .\PRDATAi[0]_4 (\PRDATAi[0]_4 ), .sercon_m_4(
        sercon_m_4), .sercon_m_0(sercon_m_0), .sercon_m_6(sercon_m_6), 
        .CoreAPB3_0_APBmslave4_PSELx(CoreAPB3_0_APBmslave4_PSELx), 
        .N_513(N_513), .N_699(N_699), .N_428(N_428), .N_529(N_529), 
        .N_411(N_411), .un12_PSELi(un12_PSELi), .un9_PRDATA_2_0(
        un9_PRDATA_2_0), .psh_enable_reg1_1_sqmuxa_0(
        psh_enable_reg1_1_sqmuxa_0), .N_629(N_629), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .N_426(N_426), .N_432(N_432), .N_685(N_685), .N_680(N_680), 
        .N_684(N_684), .N_681(N_681), .N_703(N_703), .N_698(N_698), 
        .N_702(N_702), .N_691(N_691), .CoreAPB3_0_APBmslave0_PSELx(
        CoreAPB3_0_APBmslave0_PSELx), .N_709(N_709), .N_679(N_679), 
        .N_678(N_678), .N_506(N_506), .N_711(N_711), .N_140(N_140), 
        .N_710(N_710), .un4_PRDATA(un4_PRDATA), .N_700(N_700), .N_687(
        N_687), .N_705(N_705), .N_688(N_688), .N_706(N_706), .N_690(
        N_690), .N_708(N_708), .N_689(N_689), .N_707(N_707), .N_686(
        N_686), .N_704(N_704), .PRDATA_regif_sn_N_20_i_1(
        PRDATA_regif_sn_N_20_i_1), .N_660(N_660));
    CFG4 #( .INIT(16'h0010) )  \iPSELS_0_a2[0]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13]), .C(N_426), .D(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        CoreAPB3_0_APBmslave0_PSELx));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h4) )  \iPSELS_0[1]  (.A(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15]), .B(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .Y(N_426));
    
endmodule


module COREI2CREAL_Z3_layer0(
       COREI2C_0_0_SDAO_i,
       COREI2C_0_0_SCLO_i,
       COREI2C_0_0_INT,
       CoreAPB3_0_APBmslave0_PADDR,
       sersta_m_0,
       serdat_m,
       CoreAPB3_0_APBmslave0_PWDATA,
       serdat_4,
       serdat_0,
       sersta_m_3,
       sercon_m_6,
       sercon_m_4,
       sercon_m_0,
       \PRDATAi[0]_0 ,
       \PRDATAi[0]_1 ,
       \PRDATAi[0]_2 ,
       \PRDATAi[0]_6 ,
       \PRDATAi[0]_4 ,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       un9_PRDATA_2_0,
       BIBUF_COREI2C_0_0_SDA_IO_Y,
       BIBUF_COREI2C_0_0_SCL_IO_Y,
       N_528,
       psh_enable_reg1_1_sqmuxa_0,
       un4_PRDATA,
       un12_PSELi,
       CoreAPB3_0_APBmslave1_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE
    );
output [0:0] COREI2C_0_0_SDAO_i;
output [0:0] COREI2C_0_0_SCLO_i;
output [0:0] COREI2C_0_0_INT;
input  [4:0] CoreAPB3_0_APBmslave0_PADDR;
output [1:1] sersta_m_0;
output [6:6] serdat_m;
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output serdat_4;
output serdat_0;
output sersta_m_3;
output sercon_m_6;
output sercon_m_4;
output sercon_m_0;
output \PRDATAi[0]_0 ;
output \PRDATAi[0]_1 ;
output \PRDATAi[0]_2 ;
output \PRDATAi[0]_6 ;
output \PRDATAi[0]_4 ;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output un9_PRDATA_2_0;
input  BIBUF_COREI2C_0_0_SDA_IO_Y;
input  BIBUF_COREI2C_0_0_SCL_IO_Y;
input  N_528;
input  psh_enable_reg1_1_sqmuxa_0;
output un4_PRDATA;
input  un12_PSELi;
input  CoreAPB3_0_APBmslave1_PSELx;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;

    wire \COREI2C_0_0_SDAO[0] , \COREI2C_0_0_SCLO[0] , 
        \fsmdet[3]_net_1 , \fsmdet_i_0[3] , SCLInt_net_1, SCLInt_i_0, 
        \SDAI_ff_reg[3]_net_1 , GND_net_1, \SDAI_ff_reg_3[3] , 
        VCC_net_1, \SCLI_ff_reg[0]_net_1 , \SCLI_ff_reg_3[0] , 
        \SCLI_ff_reg[1]_net_1 , \SCLI_ff_reg_3[1] , 
        \SCLI_ff_reg[2]_net_1 , \SCLI_ff_reg_3[2] , 
        \SCLI_ff_reg[3]_net_1 , \SCLI_ff_reg_3[3] , 
        \SDAI_ff_reg[0]_net_1 , \SDAI_ff_reg_3[0] , 
        \SDAI_ff_reg[1]_net_1 , \SDAI_ff_reg_3[1] , 
        \SDAI_ff_reg[2]_net_1 , \SDAI_ff_reg_3[2] , \sercon[7]_net_1 , 
        sercon18, \PCLK_count2[0]_net_1 , \PCLK_count2_4[0]_net_1 , 
        \PCLK_count2[1]_net_1 , \PCLK_count2_4[1]_net_1 , 
        \framesync[0]_net_1 , \framesync_6[0] , \framesync[1]_net_1 , 
        \framesync_6[1] , \framesync[2]_net_1 , \framesync_6[2] , 
        \framesync[3]_net_1 , \framesync_6[3] , \PCLK_count1[0]_net_1 , 
        \PCLK_count1_4[0] , \PCLK_count1[1]_net_1 , \PCLK_count1_4[1] , 
        \PCLK_count1[2]_net_1 , \PCLK_count1_4[2] , 
        \PCLK_count1[3]_net_1 , \PCLK_count1_4[3] , \indelay[0]_net_1 , 
        \indelay_4[0]_net_1 , \indelay[1]_net_1 , \indelay_4[1]_net_1 , 
        \indelay[2]_net_1 , \indelay_4[2]_net_1 , \sercon[0]_net_1 , 
        \sercon[1]_net_1 , \sercon[2]_net_1 , \sercon_9[3] , 
        \sercon[4]_net_1 , \sercon_9[4] , \sercon[5]_net_1 , 
        \sercon[6]_net_1 , \serdat[1]_net_1 , \serdat_19[1] , 
        un1_serdat_2_sqmuxa_net_1, \serdat[2]_net_1 , \serdat_19[2] , 
        \serdat[3]_net_1 , \serdat_19[3] , \serdat_19[4] , 
        \serdat[5]_net_1 , \serdat_19[5] , \serdat[6]_net_1 , 
        \serdat_19[6] , \serdat[7]_net_1 , \serdat_19[7] , 
        \serdat_19[0] , \sersta[4]_net_1 , \sersta_3[4] , sclscl_net_1, 
        \fsmmod[5]_net_1 , sclscl_1_sqmuxa_i_0, SDAInt_net_1, 
        un1_SDAInt5, un1_SCLInt5, nedetect_net_1, 
        nedetect_0_sqmuxa_net_1, SCLInt6, starto_en_net_1, starto_en8, 
        starto_en_1_sqmuxa_i_0, pedetect_net_1, 
        pedetect_0_sqmuxa_net_1, un1_SCLI_ff_reg, \fsmsta[0]_net_1 , 
        \fsmsta_9[0] , un1_ens1_pre_1_sqmuxa_i_0, \fsmsta[1]_net_1 , 
        N_1328_i_0, \fsmsta[2]_net_1 , \fsmsta_9[2] , 
        \fsmsta[3]_net_1 , N_1306_i_0, \fsmsta[4]_net_1 , 
        \fsmsta_9[4] , \sersta[0]_net_1 , \sersta_3[0] , 
        \sersta[1]_net_1 , \sersta_3[1] , \sersta[2]_net_1 , 
        \sersta_3[2] , \sersta[3]_net_1 , \sersta_3[3] , ack_net_1, 
        ack_10, N_1272, SDAO_int_1_sqmuxa_i_0, bsd7_net_1, 
        bsd7_10_iv_i_0, bsd7_tmp_net_1, bsd7_tmp_7, adrcomp_net_1, 
        un1_adrcomp14_1_net_1, adrcomp_2_sqmuxa_i_0, ack_bit_net_1, 
        ack_bit_1_sqmuxa_net_1, PCLKint_net_1, PCLKint_4, 
        un1_fsmdet_1_i_0, busfree_net_1, un1_fsmdet, adrcompen_net_1, 
        un1_adrcomp14_net_1, adrcompen_2_sqmuxa_i_0, \fsmdet[0]_net_1 , 
        \fsmdet[1]_net_1 , N_871_i_0, \fsmdet[2]_net_1 , N_873_i_0, 
        N_875_i_0, \fsmdet[4]_net_1 , N_877_i_0, \fsmdet[5]_net_1 , 
        N_879_i_0, \fsmdet[6]_net_1 , N_881_i_0, \fsmsync[0]_net_1 , 
        \fsmsync_ns[0] , \fsmsync[1]_net_1 , N_955_i_0, 
        \fsmsync[2]_net_1 , N_957_i_0, \fsmsync[3]_net_1 , N_959_i_0, 
        \fsmsync[4]_net_1 , N_961_i_0, \fsmsync[5]_net_1 , N_963_i_0, 
        \fsmsync[6]_net_1 , N_965_i_0, \fsmmod[0]_net_1 , 
        \fsmmod_ns[0] , \fsmmod[1]_net_1 , \fsmmod_ns[1] , 
        \fsmmod[2]_net_1 , N_1010_i_0, \fsmmod[3]_net_1 , 
        \fsmmod_ns[3] , \fsmmod[4]_net_1 , N_1013_i_0, \fsmmod_ns[5] , 
        \fsmmod[6]_net_1 , N_1016_i_0, PCLK_count1_ov_net_1, 
        PCLK_count1_ov_3, PCLKint_ff_net_1, PCLKint_ff_3, 
        PCLK_count2_ov_net_1, PCLK_count2_ov_0_sqmuxa_net_1, 
        SCLO_int5_i_0, framesync24, un1_sersta69_net_1, 
        un1_fsmsta_nxt_2_sn_N_3, N_756, \NoName_cnst_2[3] , 
        \un1_fsmsta_nxt_2_bm[3]_net_1 , un1_sersta58_1, 
        un1_serdat_2_sqmuxa_1_0_1_net_1, un1_sersta60_1_net_1, 
        un1_serdat_2_sqmuxa_1_1_net_1, CO1, counter_PRESETN, 
        PCLK_count17, un1_framesync24, fsmsta13, un1_adrcomp, 
        un1_PRDATA_1, \sercon_m[3] , un1_fsmmod_1, N_980, 
        counter_PRESETN_1_net_1, fsmsta_9_2_342_i_a4_0, 
        \PRDATA_0_iv_RNO_1[7]_net_1 , un14_PRDATA_net_1, 
        \PRDATA_0_iv_0[7] , un1_PRDATA, un1_sersta58, bsd7_10_iv_1, 
        bsd7_10_iv_i_1, \PWDATA_i_m_0[7] , 
        \un1_bsd7_1_sqmuxa[0]_net_1 , serdat4, 
        serdat_2_sqmuxa_1_0_net_1, fsmsta_9_2_342_i_1_1, 
        un1_sersta84_2_0, N_1306_i_1, fsmsta_9_2_342_i_a2, 
        un1_fsmsta_nxt_1_sqmuxa_net_1, N_1123, fsmsta_9_2_342_i_a2_0, 
        fsmsta_9_2_342_i_a1_1, un1_sersta65_1, sercon7_1, 
        un1_fsmmod_2_2, sercon7, fsmmod_nxt_0_sqmuxa, un1_framesync_4, 
        \un1_fsmsta_nxt_0_1_iv_1_0[2]_net_1 , 
        \un1_fsmsta_nxt_0_1_iv_1[2]_net_1 , sersta71, 
        un1_sersta60_net_1, \un1_fsmsta_nxt[2] , sersta84_2, sersta65, 
        un1_fsmsta, \sersta_3_1[3] , N_1237_2, N_1020_1, 
        un1_fsmsta_nxt_1_sqmuxa_1_1_net_1, fsmsta_nxt19, 
        un1_fsmsta_nxt_1_sqmuxa_1_net_1, fsmsta_nxt_1_sqmuxa_4_0_net_1, 
        \un1_fsmsta_nxt_2_ns_1[4]_net_1 , un1_framesync24_1_net_1, 
        N_1124, N_5, un1_sersta71_net_1, bsd7_tmp_7_am, 
        bsd7_tmp_7_ns_1, un1_fsmdet_2, \fsmsta_9_am[2] , 
        \fsmsta_9_bm[2] , \fsmsta_9_am[4] , \fsmsta_9_bm[4] , 
        framesync_6_e2, \framesync_6_enl_am[0] , 
        \framesync_6_enl_bm[0] , \framesync_6_enl_bm[3] , 
        \framesync_6_enl_am[3] , \un1_fsmsta_nxt_2_am[3]_net_1 , 
        \fsmsta_nxt_3_0_d_am[1]_net_1 , \fsmsta_nxt_3_0_d_bm[1]_net_1 , 
        \fsmsta_nxt_3_0_d_ns[1]_net_1 , N_1149, \un1_fsmsta_nxt_2[0] , 
        N_1126, N_1122, N_1151, N_1128, \fsmsta_nxt_3[0]_net_1 , 
        N_1066, un1_framesync_2, CO0, \un1_fsmsta_nxt_0_1_iv[3]_net_1 , 
        un1_sersta84_1_1_0_net_1, un1_sersta84_1_2_net_1, 
        \un1_fsmsta_nxt_1[3]_net_1 , N_827, counter_PRESETN_1_0_net_1, 
        adrcomp12, bsd7_tmp_7_sn_m6_1_0, 
        \fsmsync_ns_0_a3_3_0[0]_net_1 , sersta75_0, 
        \fsmmod_ns_i_a4_0[2] , un9_PRDATA_1_net_1, N_1236_2, 
        sersta80_1, N_1236_1, mst, PCLKint_p1_net_1, sersta77_2, 
        un14_PRDATA_2, N_1290_2, N_1059, bsd7_tmp_i_m_1, N_974, 
        N_1237_1, sersta85_1, sersta74_2, SDAO_int_6_0_312_1, 
        SDAO_int_1_sqmuxa_1_net_1, un1_fsmsync_2, un1_sercon_1_4, 
        un1_sercon_1_3, \fsmmod_ns_0_a4_0_4_0[3]_net_1 , 
        \fsmsta_cnst_i_0[4]_net_1 , \fsmsync_ns_0_a3_0_2[0]_net_1 , 
        fsmsta19_2_0, fsmsta_nxt_1_sqmuxa_5_1, 
        fsmsta_nxt_1_sqmuxa_0_net_1, sersta65_1, sersta81_0, N_1020, 
        un1_framesync_1, fsmsta33, N_1235, un18_counter_PRESETN_net_1, 
        sersta66, framesync_6_sm0, N_1023, N_1237, N_1029, N_1290_1, 
        sersta78_3, sersta77_3, N_4, N_1236, N_4_0, N_1034, 
        SDAO_int_1_sqmuxa_2_net_1, un1_sersta84_2_1_0_net_1, 
        un1_fsmdet_1_3_net_1, un1_fsmdet_1_2_net_1, 
        \fsmmod_ns_i_a4_2[2]_net_1 , \fsmmod_ns_i_a4_1[2]_net_1 , 
        \sercon_8_1[4] , \sersta_m[0] , sersta72, sersta64, sersta61, 
        fsmsta19, N_989, N_1225, N_1031, N_1052, N_999, sersta82, 
        sersta83, sersta81, sersta85, \fsmsta_nxt_4_m[2] , sersta76, 
        sersta70, sersta75, sersta74, sersta67, N_985, un1_sersta64_0, 
        sersta84, sersta69, un1_fsmdet_2_0, N_994, un1_framesync24_1_0, 
        sersta77, \fsmsta_nxt_4_i_m[0] , \fsmsta_nxt_4_i_m[3] , 
        un1_fsmdet_0, un1_fsmsta33, N_7, N_22, fsmsta_9_2_342_i_a1_0, 
        SDAO_int_1_sqmuxa_4_net_1, un1_fsmsta_nxt_1_sqmuxa_0_net_1, 
        un1_sersta65_1_0, \fsmmod_ns_i_0[4]_net_1 , 
        \fsmmod_ns_0_0[0]_net_1 , \fsmmod_ns_i_0_0[2]_net_1 , 
        \fsmsync_ns_i_0[6]_net_1 , \un1_fsmsta_nxt_0_1_iv_1[1]_net_1 , 
        fsmsta_9_2_342_i_a3_0, un1_sercon_1_6, 
        \fsmsync_ns_i_0[3]_net_1 , un1_sersta69_0, framesync10, N_972, 
        N_1224, N_990, un1_PSEL, \fsmmod_ns_0_a4_0_4[3]_net_1 , N_1049, 
        N_25_mux, un1_sersta78, \sercon_m[2] , \sersta_m[4] , 
        \sercon_m[5] , \sersta_m[2] , un1_sersta65_1_1, 
        fsmsta_nxt_1_sqmuxa_2_net_1, N_26_mux, fsmsta_nxt93, N_973, 
        N_1072, N_1223, \fsmsta_cnst_i_0[0]_net_1 , un1_sersta65_1_1_0, 
        \fsmsync_ns_i_1[6]_net_1 , fsmsta_3_sqmuxa_0_net_1, 
        \fsmsync_ns_0_1[0]_net_1 , un1_sersta64_4, un1_sersta64_3, 
        fsmmod5, N_983, un1_fsmsta_nxt_1_sqmuxa_4_net_1, un1_sercon_1, 
        fsmsta_9_2_342_i_a3, \un1_fsmsta_nxt[1] , N_1047, N_1040, 
        N_1311, CO1_0, N_1048_2, framesync14, 
        PCLK_count1_0_sqmuxa_net_1, un1_framesync24_0, 
        fsmsta_9_0_372_i_0, bsd7_tmp_i_m_1_0, N_1288, 
        \un1_fsmsta_nxt_0_0_iv[0]_net_1 , N_1110, N_6, 
        \un1_fsmsta_nxt_1[1]_net_1 , \serdat_i_m_0[7] , serdat48, 
        serdat_0_sqmuxa_net_1, adrcomp7, N_1289, 
        \un1_fsmsta_nxt_1[2]_net_1 , \un1_fsmsta_nxt_1[0]_net_1 , 
        fsmsta_9_0_372_i_m4_d, un1_serdat_2_sqmuxa_1_tz_net_1, 
        fsmsta_9_0_372_i_m4_s, fsmsta_9_0_372_i_m4_0_d, 
        un1_serdat_2_sqmuxa_1_net_1, N_1330;
    
    CFG3 #( .INIT(8'hAC) )  \un1_fsmsta_nxt_2_ns[3]  (.A(
        \un1_fsmsta_nxt_2_bm[3]_net_1 ), .B(
        \un1_fsmsta_nxt_2_am[3]_net_1 ), .C(un1_fsmsta_nxt_2_sn_N_3), 
        .Y(N_1123));
    CFG2 #( .INIT(4'hD) )  \SMBint_filter_proc.SCLI_ff_reg_3[1]  (.A(
        \sercon[6]_net_1 ), .B(\SCLI_ff_reg[0]_net_1 ), .Y(
        \SCLI_ff_reg_3[1] ));
    CFG4 #( .INIT(16'h8807) )  \un1_bsd7_1_sqmuxa[0]  (.A(un4_PRDATA), 
        .B(un1_PSEL), .C(nedetect_net_1), .D(COREI2C_0_0_INT[0]), .Y(
        \un1_bsd7_1_sqmuxa[0]_net_1 ));
    CFG2 #( .INIT(4'hB) )  \PCLKint_write_proc.PCLKint_4  (.A(
        counter_PRESETN), .B(PCLKint_net_1), .Y(PCLKint_4));
    CFG4 #( .INIT(16'h0004) )  un1_serdat_2_sqmuxa_1_1 (.A(
        un1_sersta58_1), .B(un1_serdat_2_sqmuxa_1_0_1_net_1), .C(
        \fsmdet[3]_net_1 ), .D(un1_sersta60_1_net_1), .Y(
        un1_serdat_2_sqmuxa_1_1_net_1));
    CFG3 #( .INIT(8'h31) )  \serdat_write_proc.bsd7_10_iv_i  (.A(
        un1_sersta58), .B(bsd7_10_iv_1), .C(bsd7_10_iv_i_1), .Y(
        bsd7_10_iv_i_0));
    CFG4 #( .INIT(16'h0100) )  \SDAO_int_write_proc.sersta75  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(sersta75_0), .Y(sersta75));
    SLE \sercon[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \sercon_write_proc.sercon18  (.A(un1_PSEL), 
        .B(un1_PRDATA), .Y(sercon18));
    CFG2 #( .INIT(4'hB) )  \fsmsync_ns_i_o3_0[2]  (.A(N_972), .B(
        SCLInt_net_1), .Y(N_983));
    SLE \fsmdet[1]  (.D(N_871_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[1]_net_1 ));
    CFG4 #( .INIT(16'h3ACA) )  
        \framesync_write_proc.framesync_6_enl[2]  (.A(
        \fsmdet[3]_net_1 ), .B(\framesync[2]_net_1 ), .C(
        framesync_6_e2), .D(CO1_0), .Y(\framesync_6[2] ));
    SLE SDAInt (.D(\SDAI_ff_reg[0]_net_1 ), .CLK(GL0_INST), .EN(
        un1_SDAInt5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        SDAInt_net_1));
    CFG4 #( .INIT(16'h45EF) )  \fsmsta_RNO_0[3]  (.A(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .B(N_1123), .C(
        fsmsta_9_2_342_i_a2_0), .D(fsmsta_9_2_342_i_a1_1), .Y(
        N_1306_i_1));
    SLE starto_en (.D(starto_en8), .CLK(GL0_INST), .EN(
        starto_en_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(starto_en_net_1));
    CFG1 #( .INIT(2'h1) )  SDAO_int_RNINGI9 (.A(\COREI2C_0_0_SDAO[0] ), 
        .Y(COREI2C_0_0_SDAO_i[0]));
    CFG4 #( .INIT(16'h2000) )  \sercon_write_proc.sersta84  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(sersta84_2), .D(
        \fsmsta[1]_net_1 ), .Y(sersta84));
    CFG4 #( .INIT(16'h3133) )  \un1_fsmsta_nxt_0_1_iv_1_0[2]  (.A(
        sersta84_2), .B(sersta65), .C(\fsmsta[1]_net_1 ), .D(
        un1_fsmsta), .Y(\un1_fsmsta_nxt_0_1_iv_1_0[2]_net_1 ));
    CFG3 #( .INIT(8'h08) )  \sersta_RNIBH1B1[1]  (.A(\sersta[1]_net_1 )
        , .B(CoreAPB3_0_APBmslave0_PADDR[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(sersta_m_0[1]));
    SLE \serdat[4]  (.D(\serdat_19[4] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(serdat_4));
    SLE \fsmsta[4]  (.D(\fsmsta_9[4] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\fsmsta[4]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \SDAO_int_write_proc.un1_sersta58  (.A(
        un1_sersta58_1), .B(un1_sersta60_1_net_1), .Y(un1_sersta58));
    SLE \SCLI_ff_reg[1]  (.D(\SCLI_ff_reg_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[1]_net_1 ));
    SLE pedetect (.D(pedetect_0_sqmuxa_net_1), .CLK(GL0_INST), .EN(
        un1_SCLI_ff_reg), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(pedetect_net_1));
    SLE \fsmmod[4]  (.D(N_1013_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[4]_net_1 ));
    CFG4 #( .INIT(16'hFEFF) )  \busfree_write_proc.un1_fsmdet  (.A(
        fsmmod_nxt_0_sqmuxa), .B(un1_fsmdet_2_0), .C(\fsmdet[3]_net_1 )
        , .D(\sercon[6]_net_1 ), .Y(un1_fsmdet));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_proc.SDAI_ff_reg_3[3]  (.A(
        \sercon[6]_net_1 ), .B(\SDAI_ff_reg[2]_net_1 ), .Y(
        \SDAI_ff_reg_3[3] ));
    CFG4 #( .INIT(16'h1113) )  un1_serdat_2_sqmuxa_1_tz (.A(
        COREI2C_0_0_INT[0]), .B(\fsmdet[3]_net_1 ), .C(un1_sersta58), 
        .D(un1_sersta65_1), .Y(un1_serdat_2_sqmuxa_1_tz_net_1));
    CFG4 #( .INIT(16'h0800) )  \fsmmod_ns_0_a4_0_4[3]  (.A(
        \fsmmod_ns_0_a4_0_4_0[3]_net_1 ), .B(N_1020), .C(N_1029), .D(
        un1_framesync_2), .Y(\fsmmod_ns_0_a4_0_4[3]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \fsmmod_ns_0[0]  (.A(N_1031), .B(
        \fsmmod[0]_net_1 ), .C(fsmmod5), .D(\fsmmod_ns_0_0[0]_net_1 ), 
        .Y(\fsmmod_ns[0] ));
    CFG4 #( .INIT(16'hECCC) )  \fsmmod_ns_0_0[0]  (.A(
        \fsmmod[5]_net_1 ), .B(fsmmod_nxt_0_sqmuxa), .C(sclscl_net_1), 
        .D(pedetect_net_1), .Y(\fsmmod_ns_0_0[0]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \SDAO_int_write_proc.sersta67  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(N_1236_2), .Y(sersta67));
    SLE ack (.D(ack_10), .CLK(GL0_INST), .EN(\sercon[6]_net_1 ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(ack_net_1));
    CFG4 #( .INIT(16'h0100) )  \adrcomp_write_proc.sersta74  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .D(N_1237_1), .Y(sersta74));
    CFG3 #( .INIT(8'hAB) )  \SDAO_int_write_proc.un1_sersta58_1  (.A(
        un1_sersta78), .B(\fsmsta[1]_net_1 ), .C(N_1020_1), .Y(
        un1_sersta58_1));
    CFG4 #( .INIT(16'h7FFF) )  \SCLInt_write_proc.SCLInt6  (.A(
        \SCLI_ff_reg[0]_net_1 ), .B(\SCLI_ff_reg[3]_net_1 ), .C(
        \SCLI_ff_reg[2]_net_1 ), .D(\SCLI_ff_reg[1]_net_1 ), .Y(
        SCLInt6));
    SLE \fsmsta[3]  (.D(N_1306_i_0), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\fsmsta[3]_net_1 ));
    CFG4 #( .INIT(16'h335F) )  \un1_fsmsta_nxt_2_ns_1[4]  (.A(
        framesync24), .B(N_5), .C(un1_sersta71_net_1), .D(
        un1_fsmsta_nxt_2_sn_N_3), .Y(\un1_fsmsta_nxt_2_ns_1[4]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \SDAO_int_write_proc.sersta60_1  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[4]_net_1 ), .Y(N_1236_1));
    CFG4 #( .INIT(16'h0E00) )  \serdat_write_proc.bsd7_10_iv_1_RNO  (
        .A(un1_sersta60_1_net_1), .B(un1_sersta58_1), .C(
        bsd7_tmp_net_1), .D(bsd7_tmp_i_m_1), .Y(bsd7_tmp_i_m_1_0));
    CFG4 #( .INIT(16'hECCC) )  \un1_fsmsta_nxt_0_1_iv_1[2]  (.A(N_1235)
        , .B(\fsmsta_nxt_4_m[2] ), .C(\fsmsta[0]_net_1 ), .D(
        \fsmsta[1]_net_1 ), .Y(\un1_fsmsta_nxt_0_1_iv_1[2]_net_1 ));
    SLE \serdat[2]  (.D(\serdat_19[2] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  un9_PRDATA_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(un9_PRDATA_1_net_1));
    CFG4 #( .INIT(16'h4C00) )  un1_serdat_2_sqmuxa_1_0_1 (.A(
        COREI2C_0_0_INT[0]), .B(pedetect_net_1), .C(un1_sersta65_1), 
        .D(\sercon[6]_net_1 ), .Y(un1_serdat_2_sqmuxa_1_0_1_net_1));
    CFG4 #( .INIT(16'h3336) )  \sercon_write_proc.un1_framesync24  (.A(
        \framesync[2]_net_1 ), .B(\framesync[3]_net_1 ), .C(
        \framesync[1]_net_1 ), .D(\framesync[0]_net_1 ), .Y(
        un1_framesync24));
    CFG2 #( .INIT(4'hE) )  \fsmsta_sync_proc.un1_fsmdet_2  (.A(
        un1_framesync24_0), .B(un1_fsmdet_0), .Y(un1_fsmdet_2));
    CFG2 #( .INIT(4'hE) )  counter_PRESETN_1 (.A(\fsmdet[3]_net_1 ), 
        .B(\fsmdet[5]_net_1 ), .Y(counter_PRESETN_1_net_1));
    CFG2 #( .INIT(4'h8) )  \fsmsync_ns_0_a3_0[0]  (.A(
        \fsmsync_ns_0_a3_0_2[0]_net_1 ), .B(N_1059), .Y(N_985));
    CFG4 #( .INIT(16'hFFFE) )  \adrcomp_write_proc.un1_sersta64_4  (.A(
        sersta82), .B(sersta77), .C(sersta74), .D(sersta64), .Y(
        un1_sersta64_4));
    CFG4 #( .INIT(16'h0400) )  fsmsta_nxt_1_sqmuxa_2 (.A(
        \fsmsta[2]_net_1 ), .B(N_1236_1), .C(fsmsta_nxt19), .D(
        sersta74_2), .Y(fsmsta_nxt_1_sqmuxa_2_net_1));
    CFG2 #( .INIT(4'h4) )  PCLK_count1_0_sqmuxa (.A(counter_PRESETN), 
        .B(PCLK_count17), .Y(PCLK_count1_0_sqmuxa_net_1));
    CFG4 #( .INIT(16'h3953) )  \sersta_write_proc.sersta_2_4_0_.m15  (
        .A(\fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(sersta84_2), 
        .D(\fsmsta[1]_net_1 ), .Y(N_26_mux));
    CFG3 #( .INIT(8'hD8) )  \fsmsta_sync_proc.fsmsta_9_am[2]  (.A(
        un1_sersta84_2_0), .B(\un1_fsmsta_nxt_1[2]_net_1 ), .C(N_1128), 
        .Y(\fsmsta_9_am[2] ));
    CFG4 #( .INIT(16'hEEEA) )  \adrcomp_write_proc.adrcomp7  (.A(
        counter_PRESETN_1_net_1), .B(COREI2C_0_0_INT[0]), .C(
        un1_sersta64_4), .D(un1_sersta64_3), .Y(adrcomp7));
    CFG4 #( .INIT(16'h1000) )  \adrcomp_write_proc.sersta83  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(sersta84_2), .D(
        \fsmsta[1]_net_1 ), .Y(sersta83));
    CFG4 #( .INIT(16'hFF02) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_0  (
        .A(counter_PRESETN_1_net_1), .B(adrcomp_net_1), .C(fsmsta13), 
        .D(un1_fsmsta33), .Y(fsmsta_9_0_372_i_0));
    CFG3 #( .INIT(8'h15) )  SDAO_int_1_sqmuxa_4 (.A(\fsmmod[1]_net_1 ), 
        .B(adrcompen_net_1), .C(adrcomp_net_1), .Y(N_1290_1));
    CFG4 #( .INIT(16'hA0B0) )  \fsmsta_sync_proc.fsmsta13  (.A(
        adrcomp_net_1), .B(\fsmmod[0]_net_1 ), .C(un1_framesync24), .D(
        \fsmmod[5]_net_1 ), .Y(fsmsta13));
    CFG4 #( .INIT(16'hFFF2) )  un1_fsmsta_nxt_1_sqmuxa (.A(sersta61), 
        .B(fsmsta_nxt19), .C(un1_fsmsta_nxt_1_sqmuxa_4_net_1), .D(
        un1_fsmsta_nxt_1_sqmuxa_1_net_1), .Y(
        un1_fsmsta_nxt_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'hFFFE) )  un1_sersta84_2_1 (.A(N_1225), .B(
        un1_sersta84_2_1_0_net_1), .C(N_1224), .D(N_1223), .Y(
        un1_sersta84_2_0));
    CFG4 #( .INIT(16'h3313) )  \fsmsta_cnst_i[0]  (.A(fsmsta13), .B(
        \fsmsta_cnst_i_0[0]_net_1 ), .C(counter_PRESETN_1_net_1), .D(
        un1_fsmsta33), .Y(N_1066));
    CFG4 #( .INIT(16'h0001) )  un14_PRDATA (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(N_528), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(un14_PRDATA_net_1));
    CFG4 #( .INIT(16'h000D) )  \fsmsync_ns_i_a3_0[2]  (.A(
        \fsmsync[2]_net_1 ), .B(PCLKint_p1_net_1), .C(
        \fsmsync[1]_net_1 ), .D(\fsmsync[0]_net_1 ), .Y(N_989));
    CFG2 #( .INIT(4'h8) )  \fsmsta_sync_proc.un1_framesync24_1  (.A(
        framesync24), .B(adrcomp_net_1), .Y(un1_framesync24_1_0));
    CFG4 #( .INIT(16'h0400) )  \SDAO_int_write_proc.un1_framesync_2  (
        .A(\framesync[2]_net_1 ), .B(\framesync[3]_net_1 ), .C(
        \framesync[1]_net_1 ), .D(\framesync[0]_net_1 ), .Y(
        un1_framesync_2));
    CFG4 #( .INIT(16'hF0EE) )  \sercon_write_proc.sercon_9[3]  (.A(
        COREI2C_0_0_INT[0]), .B(sercon7), .C(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .D(sercon18), .Y(
        \sercon_9[3] ));
    CFG3 #( .INIT(8'hE4) )  \fsmsta_sync_proc.fsmsta_9_ns[4]  (.A(
        un1_fsmdet_2), .B(\fsmsta_9_am[4] ), .C(\fsmsta_9_bm[4] ), .Y(
        \fsmsta_9[4] ));
    SLE \fsmmod[3]  (.D(\fsmmod_ns[3] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[3]_net_1 ));
    CFG4 #( .INIT(16'hAEFF) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_o4_0  (.A(bsd7_net_1), 
        .B(\framesync[3]_net_1 ), .C(un1_framesync_2), .D(un1_sersta58)
        , .Y(N_1288));
    CFG4 #( .INIT(16'h0105) )  \framesync_write_proc.framesync_6_e2  (
        .A(un1_framesync_2), .B(nedetect_net_1), .C(framesync_6_sm0), 
        .D(framesync24), .Y(framesync_6_e2));
    CFG4 #( .INIT(16'h8000) )  \adrcomp_write_proc.un1_sercon_1_3  (.A(
        \serdat[6]_net_1 ), .B(\serdat[1]_net_1 ), .C(
        \sercon[2]_net_1 ), .D(adrcompen_net_1), .Y(un1_sercon_1_3));
    CFG4 #( .INIT(16'h1000) )  \adrcomp_write_proc.un1_sercon_1_6  (.A(
        serdat_0), .B(\serdat[2]_net_1 ), .C(un1_sercon_1_4), .D(
        un1_sercon_1_3), .Y(un1_sercon_1_6));
    CFG2 #( .INIT(4'h4) )  \sersta_write_proc.sersta85_2  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[4]_net_1 ), .Y(N_1237_1));
    CFG2 #( .INIT(4'h2) )  \SDAO_int_write_proc.sersta80_2  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(sersta77_2));
    CFG3 #( .INIT(8'h02) )  \un1_fsmsta_nxt_0_1_iv_1_RNO[2]  (.A(
        ack_net_1), .B(SDAInt_net_1), .C(N_1020), .Y(
        \fsmsta_nxt_4_m[2] ));
    CFG4 #( .INIT(16'h737F) )  \sersta_write_proc.sersta_3_1[3]  (.A(
        N_1237_2), .B(\fsmsta[1]_net_1 ), .C(sersta84_2), .D(
        un1_fsmsta), .Y(\sersta_3_1[3] ));
    CFG3 #( .INIT(8'h4E) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_m4  (.A(
        fsmsta_9_0_372_i_m4_s), .B(fsmsta_9_0_372_i_m4_d), .C(
        fsmsta_9_0_372_i_m4_0_d), .Y(N_1330));
    SLE \serdat[7]  (.D(\serdat_19[7] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[7]_net_1 ));
    CFG4 #( .INIT(16'hCC08) )  un1_fsmsta_nxt_1_sqmuxa_0 (.A(
        un1_fsmsta), .B(fsmsta_nxt_1_sqmuxa_5_1), .C(\fsmsta[3]_net_1 )
        , .D(fsmsta_nxt_1_sqmuxa_0_net_1), .Y(
        un1_fsmsta_nxt_1_sqmuxa_0_net_1));
    SLE \sercon[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[2]_net_1 ));
    CFG4 #( .INIT(16'hCCC4) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_a1_0  (.A(framesync24), .B(
        fsmsta_9_2_342_i_a4_0), .C(\sercon[2]_net_1 ), .D(SDAInt_net_1)
        , .Y(fsmsta_9_2_342_i_a1_0));
    CFG4 #( .INIT(16'hF0F8) )  counter_PRESETN_1_0 (.A(
        \fsmmod[4]_net_1 ), .B(\COREI2C_0_0_SCLO[0] ), .C(
        un18_counter_PRESETN_net_1), .D(SCLInt_net_1), .Y(
        counter_PRESETN_1_0_net_1));
    CFG2 #( .INIT(4'h8) )  \SDAO_int_write_proc.sersta63_1  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .Y(un1_fsmsta));
    CFG4 #( .INIT(16'hC400) )  \adrcomp_write_proc.un1_sercon_1_8  (.A(
        mst), .B(un1_framesync_1), .C(sersta64), .D(un1_sercon_1_6), 
        .Y(un1_sercon_1));
    CFG3 #( .INIT(8'hCA) )  \fsmsta_RNO[0]  (.A(
        \fsmsta_nxt_3[0]_net_1 ), .B(N_1066), .C(un1_fsmdet_2), .Y(
        \fsmsta_9[0] ));
    CFG4 #( .INIT(16'h1101) )  fsmsta_nxt_1_sqmuxa_1_0 (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(
        \COREI2C_0_0_SDAO[0] ), .D(SDAInt_net_1), .Y(
        fsmsta_nxt_1_sqmuxa_5_1));
    CFG3 #( .INIT(8'h40) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_a2  (.A(
        \un1_fsmsta_nxt_1[3]_net_1 ), .B(fsmsta_9_2_342_i_a2_0), .C(
        un1_sersta84_2_0), .Y(fsmsta_9_2_342_i_a2));
    CFG4 #( .INIT(16'h0600) )  \PCLK_counter1_proc.PCLK_count1_4[1]  (
        .A(\PCLK_count1[0]_net_1 ), .B(\PCLK_count1[1]_net_1 ), .C(
        counter_PRESETN), .D(PCLK_count17), .Y(\PCLK_count1_4[1] ));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_proc.SDAI_ff_reg_3[2]  (.A(
        \sercon[6]_net_1 ), .B(\SDAI_ff_reg[1]_net_1 ), .Y(
        \SDAI_ff_reg_3[2] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h04) )  \serdat_write_proc.serdat48  (.A(
        \fsmdet[3]_net_1 ), .B(un1_sersta65_1), .C(un1_sersta58), .Y(
        serdat48));
    CFG3 #( .INIT(8'h80) )  \fsmsta_comb_proc.fsmsta_nxt93  (.A(
        adrcompen_net_1), .B(adrcomp_net_1), .C(framesync24), .Y(
        fsmsta_nxt93));
    CFG4 #( .INIT(16'h0080) )  \PRDATA_0_iv_RNO[3]  (.A(
        un9_PRDATA_1_net_1), .B(un9_PRDATA_2_0), .C(\sersta[0]_net_1 ), 
        .D(CoreAPB3_0_APBmslave0_PADDR[0]), .Y(\sersta_m[0] ));
    CFG4 #( .INIT(16'hCCD8) )  \fsmsta_sync_proc.fsmsta_9_am[4]  (.A(
        un1_sersta84_2_0), .B(\fsmsta[4]_net_1 ), .C(N_1124), .D(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .Y(\fsmsta_9_am[4] ));
    SLE sclscl (.D(\fsmmod[5]_net_1 ), .CLK(GL0_INST), .EN(
        sclscl_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sclscl_net_1));
    CFG4 #( .INIT(16'hFF40) )  \fsmmod_ns_i_0[4]  (.A(
        \fsmmod[2]_net_1 ), .B(SCLInt_net_1), .C(PCLKint_p1_net_1), .D(
        N_1034), .Y(\fsmmod_ns_i_0[4]_net_1 ));
    CFG3 #( .INIT(8'h12) )  \PCLK_count2_4[0]  (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN), .C(
        \PCLK_count2[0]_net_1 ), .Y(\PCLK_count2_4[0]_net_1 ));
    CFG4 #( .INIT(16'h0015) )  \framesync_write_proc.framesync10  (.A(
        COREI2C_0_0_INT[0]), .B(N_1020), .C(\sercon[5]_net_1 ), .D(
        \sercon[4]_net_1 ), .Y(framesync10));
    CFG1 #( .INIT(2'h1) )  busfree_RNO (.A(\fsmdet[3]_net_1 ), .Y(
        \fsmdet_i_0[3] ));
    CFG2 #( .INIT(4'h1) )  un1_adrcomp14_1 (.A(adrcomp7), .B(adrcomp12)
        , .Y(un1_adrcomp14_1_net_1));
    SLE \SCLI_ff_reg[0]  (.D(\SCLI_ff_reg_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \fsmsync_sync_proc.un1_sersta69_1_a5_1  
        (.A(\fsmsta[3]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .D(\fsmsta[1]_net_1 ), .Y(N_1236));
    CFG4 #( .INIT(16'h00AE) )  \fsmsync_RNO[6]  (.A(\fsmsync[6]_net_1 )
        , .B(\sercon[4]_net_1 ), .C(N_973), .D(
        \fsmsync_ns_i_1[6]_net_1 ), .Y(N_965_i_0));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_proc.SDAI_ff_reg_3[0]  (.A(
        \sercon[6]_net_1 ), .B(BIBUF_COREI2C_0_0_SDA_IO_Y), .Y(
        \SDAI_ff_reg_3[0] ));
    CFG4 #( .INIT(16'hAA8A) )  \sercon_write_proc.sercon7  (.A(
        \sercon[6]_net_1 ), .B(un1_fsmmod_1), .C(sercon7_1), .D(
        un1_fsmmod_2_2), .Y(sercon7));
    CFG3 #( .INIT(8'h51) )  \fsmmod_ns_i_a4[6]  (.A(\fsmmod[6]_net_1 ), 
        .B(\fsmmod[3]_net_1 ), .C(N_1023), .Y(N_1049));
    CFG4 #( .INIT(16'hFFFD) )  counter_PRESETN_1_0_RNIIM8F (.A(N_827), 
        .B(counter_PRESETN_1_net_1), .C(counter_PRESETN_1_0_net_1), .D(
        adrcomp12), .Y(counter_PRESETN));
    CFG2 #( .INIT(4'hE) )  \fsmmod_ns_i_o4_1_1[2]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_1020_1));
    SLE \SCLI_ff_reg[3]  (.D(\SCLI_ff_reg_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[3]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  SDAO_int_1_sqmuxa_i (.A(
        SDAO_int_1_sqmuxa_1_net_1), .B(SDAO_int_1_sqmuxa_2_net_1), .C(
        SDAO_int_1_sqmuxa_4_net_1), .D(un1_sersta65_1), .Y(
        SDAO_int_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'h1333) )  \sercon_write_proc.sercon7_1  (.A(
        counter_PRESETN_1_net_1), .B(fsmmod_nxt_0_sqmuxa), .C(
        adrcomp_net_1), .D(un1_framesync_4), .Y(sercon7_1));
    CFG4 #( .INIT(16'hFFFE) )  \fsmsync_sync_proc.un1_fsmsync_2  (.A(
        \fsmsync[5]_net_1 ), .B(\fsmsync[2]_net_1 ), .C(
        \fsmsync[1]_net_1 ), .D(\fsmsync[6]_net_1 ), .Y(un1_fsmsync_2));
    CFG4 #( .INIT(16'h0001) )  \fsmsync_ns_0_a3_0_2[0]  (.A(
        \fsmmod[2]_net_1 ), .B(\fsmmod[3]_net_1 ), .C(
        \fsmmod[5]_net_1 ), .D(\fsmmod[4]_net_1 ), .Y(
        \fsmsync_ns_0_a3_0_2[0]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \fsmmod_ns_i_a3_0[2]  (.A(
        \sercon[4]_net_1 ), .B(COREI2C_0_0_INT[0]), .C(N_1059), .D(
        un1_framesync_2), .Y(N_1052));
    CFG2 #( .INIT(4'h8) )  \fsmmod_ns_0_a4_0_4_1[3]  (.A(
        \fsmmod_ns_i_a4_0[2] ), .B(\fsmmod[2]_net_1 ), .Y(
        \fsmmod_ns_0_a4_0_4_0[3]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \adrcomp_write_proc.sersta82_0  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .Y(N_1237_2));
    CFG3 #( .INIT(8'hDF) )  PCLKint_RNO (.A(un1_fsmdet_1_3_net_1), .B(
        adrcomp12), .C(un1_fsmdet_1_2_net_1), .Y(un1_fsmdet_1_i_0));
    CFG3 #( .INIT(8'h40) )  PCLKint_ff_RNIPEFR (.A(PCLKint_net_1), .B(
        \fsmmod[4]_net_1 ), .C(PCLKint_ff_net_1), .Y(fsmsta33));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[5]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .B(serdat_4), .C(un1_PSEL), 
        .D(un4_PRDATA), .Y(\serdat_19[5] ));
    CFG4 #( .INIT(16'h2000) )  \SDAO_int_write_proc.un1_framesync_1  (
        .A(\framesync[2]_net_1 ), .B(\framesync[3]_net_1 ), .C(
        \framesync[1]_net_1 ), .D(\framesync[0]_net_1 ), .Y(
        un1_framesync_1));
    CFG3 #( .INIT(8'h07) )  \fsmmod_ns_i_o4_1_RNIEV1Q[2]  (.A(
        ack_net_1), .B(SDAInt_net_1), .C(N_1020), .Y(
        \fsmsta_nxt_4_i_m[3] ));
    CFG2 #( .INIT(4'h8) )  \PCLK_count1_RNI3ADA[1]  (.A(
        \PCLK_count1[0]_net_1 ), .B(\PCLK_count1[1]_net_1 ), .Y(CO1));
    CFG4 #( .INIT(16'hEEE2) )  \fsmsta_nxt_3_0_d_bm[1]  (.A(
        \fsmsta[1]_net_1 ), .B(framesync24), .C(\sercon[2]_net_1 ), .D(
        SDAInt_net_1), .Y(\fsmsta_nxt_3_0_d_bm[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \sercon_write_proc.adrcomp12  (.A(mst), .B(
        \sercon[4]_net_1 ), .Y(adrcomp12));
    CFG4 #( .INIT(16'hFFEA) )  un1_fsmsta_nxt_1_sqmuxa_4 (.A(
        fsmsta_nxt_1_sqmuxa_2_net_1), .B(framesync24), .C(un1_sersta78)
        , .D(un1_fsmsta_nxt_1_sqmuxa_0_net_1), .Y(
        un1_fsmsta_nxt_1_sqmuxa_4_net_1));
    CFG3 #( .INIT(8'h51) )  \fsmsta_RNO[1]  (.A(fsmsta_9_0_372_i_0), 
        .B(N_1330), .C(counter_PRESETN_1_net_1), .Y(N_1328_i_0));
    CFG2 #( .INIT(4'h8) )  \serdat_write_proc.serdat4  (.A(un1_PSEL), 
        .B(un4_PRDATA), .Y(serdat4));
    SLE \PCLK_count2[0]  (.D(\PCLK_count2_4[0]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\PCLK_count2[0]_net_1 ));
    SLE \sersta[0]  (.D(\sersta_3[0] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[0]_net_1 ));
    CFG4 #( .INIT(16'h7F40) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_m5  (.A(ack_bit_net_1), 
        .B(un1_framesync_1), .C(un1_sersta65_1), .D(N_1288), .Y(N_1289)
        );
    SLE \PCLK_count1[3]  (.D(\PCLK_count1_4[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[3]_net_1 ));
    SLE \indelay[2]  (.D(\indelay_4[2]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[2]_net_1 ));
    SLE \fsmsync[2]  (.D(N_957_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[2]_net_1 ));
    CFG4 #( .INIT(16'h3777) )  \fsmsync_sync_proc.SCLO_int5_i  (.A(
        un1_fsmsync_2), .B(\sercon[6]_net_1 ), .C(un1_sersta69_0), .D(
        bsd7_tmp_i_m_1), .Y(SCLO_int5_i_0));
    CFG3 #( .INIT(8'h80) )  \sercon_write_proc.un1_PRDATA_1_RNI10RD  (
        .A(un1_PRDATA_1), .B(\sercon[6]_net_1 ), .C(un14_PRDATA_2), .Y(
        sercon_m_6));
    CFG4 #( .INIT(16'hE000) )  \fsmdet_RNO[5]  (.A(\fsmdet[2]_net_1 ), 
        .B(\fsmdet[4]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_879_i_0));
    CFG4 #( .INIT(16'hFFFE) )  \framesync_write_proc.framesync14  (.A(
        sersta77_3), .B(sersta82), .C(sersta74), .D(sersta76), .Y(
        framesync14));
    SLE \framesync[3]  (.D(\framesync_6[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[3]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \SMBint_filter_proc.SCLI_ff_reg_3[0]  (.A(
        \sercon[6]_net_1 ), .B(BIBUF_COREI2C_0_0_SCL_IO_Y), .Y(
        \SCLI_ff_reg_3[0] ));
    CFG4 #( .INIT(16'hFF80) )  \un1_fsmsta_nxt_0_1_iv_1[1]  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(N_1235), .D(
        sersta83), .Y(\un1_fsmsta_nxt_0_1_iv_1[1]_net_1 ));
    CFG4 #( .INIT(16'hEB41) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_m4_d  (.A(un1_framesync24_0)
        , .B(un1_fsmsta_nxt_2_sn_N_3), .C(\COREI2C_0_0_SDAO[0] ), .D(
        N_1072), .Y(fsmsta_9_0_372_i_m4_d));
    CFG4 #( .INIT(16'h7F2A) )  \un1_fsmsta_nxt_2[2]  (.A(
        un1_fsmsta_nxt_2_sn_N_3), .B(un1_framesync24_1_net_1), .C(
        \COREI2C_0_0_SDAO[0] ), .D(N_1110), .Y(N_1122));
    CFG4 #( .INIT(16'hCCD8) )  \un1_fsmsta_nxt_1[1]  (.A(
        un1_sersta84_1_1_0_net_1), .B(\fsmsta[1]_net_1 ), .C(
        \un1_fsmsta_nxt[1] ), .D(un1_sersta84_1_2_net_1), .Y(
        \un1_fsmsta_nxt_1[1]_net_1 ));
    CFG4 #( .INIT(16'hF870) )  \serdat_write_proc.serdat_19[0]  (.A(
        un4_PRDATA), .B(un1_PSEL), .C(ack_net_1), .D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .Y(\serdat_19[0] ));
    CFG3 #( .INIT(8'h20) )  \un1_framesync_1_1.CO0  (.A(nedetect_net_1)
        , .B(un1_framesync_2), .C(\framesync[0]_net_1 ), .Y(CO0));
    CFG2 #( .INIT(4'h7) )  \fsmsync_ns_i_o3_1[3]  (.A(
        \indelay[1]_net_1 ), .B(\indelay[2]_net_1 ), .Y(N_974));
    CFG4 #( .INIT(16'hF700) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_a1_1  (.A(adrcompen_net_1), 
        .B(un1_framesync24_1_0), .C(sersta64), .D(
        fsmsta_9_2_342_i_a1_0), .Y(fsmsta_9_2_342_i_a1_1));
    CFG2 #( .INIT(4'h8) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_a3_0  (
        .A(fsmsta_9_2_342_i_a4_0), .B(ack_net_1), .Y(
        fsmsta_9_2_342_i_a3_0));
    SLE PCLK_count1_ov (.D(PCLK_count1_ov_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PCLK_count1_ov_net_1));
    CFG3 #( .INIT(8'hB8) )  \fsmsta_sync_proc.fsmsta_9_0_372_i_m4_0_d  
        (.A(\un1_fsmsta_nxt_1[1]_net_1 ), .B(un1_sersta84_2_0), .C(
        \fsmsta_nxt_3_0_d_ns[1]_net_1 ), .Y(fsmsta_9_0_372_i_m4_0_d));
    SLE \indelay[1]  (.D(\indelay_4[1]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[1]_net_1 ));
    CFG3 #( .INIT(8'hA2) )  \NoName_cnst_2_4_3__NoName_cnst_2_1_0_.m3  
        (.A(\fsmsta[4]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(
        SDAInt_net_1), .Y(N_4));
    CFG3 #( .INIT(8'hF2) )  \fsmsync_ns_i_0[6]  (.A(\fsmsync[6]_net_1 )
        , .B(SDAInt_net_1), .C(N_985), .Y(\fsmsync_ns_i_0[6]_net_1 ));
    SLE \serdat[0]  (.D(\serdat_19[0] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(serdat_0));
    CFG4 #( .INIT(16'hCE0A) )  \fsmsta_cnst_i_0[0]  (.A(ack_net_1), .B(
        \fsmmod[1]_net_1 ), .C(un1_fsmdet_0), .D(\fsmdet[3]_net_1 ), 
        .Y(\fsmsta_cnst_i_0[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \SDAO_int_write_proc.sersta67_1  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(N_1236_2));
    CFG2 #( .INIT(4'h1) )  \fsmmod_ns_i_a2[2]  (.A(\fsmmod[1]_net_1 ), 
        .B(\fsmmod[6]_net_1 ), .Y(N_1059));
    CFG3 #( .INIT(8'hB7) )  \fsmmod_ns_0_o4[3]  (.A(PCLKint_net_1), .B(
        SCLInt_net_1), .C(PCLKint_ff_net_1), .Y(N_1023));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv[1]  (.A(\sercon[1]_net_1 ), 
        .B(\serdat[1]_net_1 ), .C(un1_PRDATA), .D(un4_PRDATA), .Y(
        \PRDATAi[0]_0 ));
    SLE \framesync[2]  (.D(\framesync_6[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[2]_net_1 ));
    CFG4 #( .INIT(16'h0700) )  \fsmmod_ns_0_a4[5]  (.A(pedetect_net_1), 
        .B(sclscl_net_1), .C(fsmmod5), .D(\fsmmod[5]_net_1 ), .Y(
        N_1047));
    CFG4 #( .INIT(16'h0F07) )  un1_fsmdet_1_3 (.A(\fsmmod[4]_net_1 ), 
        .B(\COREI2C_0_0_SCLO[0] ), .C(un18_counter_PRESETN_net_1), .D(
        SCLInt_net_1), .Y(un1_fsmdet_1_3_net_1));
    CFG4 #( .INIT(16'hFF40) )  \SDAO_int_write_proc.un1_sersta78  (.A(
        \fsmsta[0]_net_1 ), .B(sersta77_2), .C(sersta80_1), .D(
        sersta78_3), .Y(un1_sersta78));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_0_iv[3]  (.A(\serdat[3]_net_1 ), 
        .B(\sersta_m[0] ), .C(\sercon_m[3] ), .D(un4_PRDATA), .Y(
        \PRDATAi[0]_2 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hAF27) )  \fsmmod_ns_i_m4[4]  (.A(
        \fsmmod[2]_net_1 ), .B(\sercon[4]_net_1 ), .C(
        \fsmmod[4]_net_1 ), .D(COREI2C_0_0_INT[0]), .Y(N_1034));
    CFG3 #( .INIT(8'h09) )  \un1_fsmsta_nxt_0_0_iv_RNO[0]  (.A(
        ack_net_1), .B(SDAInt_net_1), .C(N_1020), .Y(
        \fsmsta_nxt_4_i_m[0] ));
    CFG4 #( .INIT(16'h8001) )  \SDAInt_write_proc.un1_SDAInt5  (.A(
        \SDAI_ff_reg[3]_net_1 ), .B(\SDAI_ff_reg[2]_net_1 ), .C(
        \SDAI_ff_reg[1]_net_1 ), .D(\SDAI_ff_reg[0]_net_1 ), .Y(
        un1_SDAInt5));
    CFG4 #( .INIT(16'h1D3F) )  
        \NoName_cnst_2_4_3__NoName_cnst_2_1_0_.m5  (.A(N_4), .B(
        fsmsta_nxt93), .C(ack_net_1), .D(\fsmsta[0]_net_1 ), .Y(N_6));
    CFG4 #( .INIT(16'hFF80) )  un1_sersta69 (.A(\fsmsta[0]_net_1 ), .B(
        \fsmsta[1]_net_1 ), .C(N_1235), .D(un1_sersta65_1_1), .Y(
        un1_sersta69_net_1));
    CFG3 #( .INIT(8'h15) )  \fsmsync_ns_i_a3[5]  (.A(
        \fsmsync[5]_net_1 ), .B(\fsmsync[2]_net_1 ), .C(
        PCLKint_p1_net_1), .Y(N_994));
    CFG3 #( .INIT(8'hFE) )  adrcomp_2_sqmuxa_i (.A(adrcomp12), .B(
        un1_sercon_1), .C(adrcomp7), .Y(adrcomp_2_sqmuxa_i_0));
    SLE \sersta[1]  (.D(\sersta_3[1] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[1]_net_1 ));
    CFG4 #( .INIT(16'h5557) )  \PCLK_counter1_proc.PCLK_count17_1.CO3  
        (.A(\PCLK_count1[3]_net_1 ), .B(\PCLK_count1[2]_net_1 ), .C(
        \PCLK_count1[1]_net_1 ), .D(\PCLK_count1[0]_net_1 ), .Y(
        PCLK_count17));
    CFG3 #( .INIT(8'hBA) )  \SDAO_int_write_proc.un1_sersta65_1_1  (.A(
        sersta70), .B(\fsmsta[2]_net_1 ), .C(N_1236), .Y(
        un1_sersta65_1_1));
    SLE \fsmdet[4]  (.D(N_877_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[4]_net_1 ));
    SLE \indelay[0]  (.D(\indelay_4[0]_net_1 ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \indelay[0]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \adrcomp_write_proc.un1_sersta64_3  (.A(
        sersta83), .B(sersta76), .C(sersta81), .Y(un1_sersta64_3));
    SLE \fsmdet[0]  (.D(SCLInt_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[0]_net_1 ));
    SLE \sercon[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[7]_net_1 ));
    CFG3 #( .INIT(8'hBA) )  \fsmsta_sync_proc.fsmsta_9_bm[2]  (.A(
        fsmsta33), .B(counter_PRESETN_1_net_1), .C(N_1072), .Y(
        \fsmsta_9_bm[2] ));
    SLE ack_bit (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), 
        .EN(ack_bit_1_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(ack_bit_net_1));
    SLE \fsmsta[2]  (.D(\fsmsta_9[2] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\fsmsta[2]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \serdat_RNIFRE11[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(\serdat[6]_net_1 ), .C(
        un9_PRDATA_2_0), .D(psh_enable_reg1_1_sqmuxa_0), .Y(
        serdat_m[6]));
    CFG4 #( .INIT(16'hF7F3) )  
        \SDAO_int_write_proc.SDAO_int_6_0_312_1  (.A(adrcomp_net_1), 
        .B(\sercon[6]_net_1 ), .C(\fsmmod[3]_net_1 ), .D(
        \fsmmod[0]_net_1 ), .Y(SDAO_int_6_0_312_1));
    SLE \fsmdet[2]  (.D(N_873_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \fsmmod_ns_0_a4_0_4_0[3]  (.A(PCLKint_net_1)
        , .B(PCLKint_ff_net_1), .Y(\fsmmod_ns_i_a4_0[2] ));
    CFG4 #( .INIT(16'h0E00) )  \fsmdet_RNO[2]  (.A(\fsmdet[0]_net_1 ), 
        .B(\fsmdet[2]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_873_i_0));
    SLE \framesync[1]  (.D(\framesync_6[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \fsmsta_sync_proc.fsmsta_9_ns[2]  (.A(
        un1_fsmdet_2), .B(\fsmsta_9_am[2] ), .C(\fsmsta_9_bm[2] ), .Y(
        \fsmsta_9[2] ));
    CFG3 #( .INIT(8'h01) )  fsmsta_nxt_1_sqmuxa_0 (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .Y(fsmsta_nxt_1_sqmuxa_0_net_1));
    CFG2 #( .INIT(4'h1) )  un9_PRDATA_2_0_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(un9_PRDATA_2_0));
    CFG4 #( .INIT(16'h0080) )  \PRDATA_0_iv_RNO[7]  (.A(
        un9_PRDATA_1_net_1), .B(un9_PRDATA_2_0), .C(\sersta[4]_net_1 ), 
        .D(CoreAPB3_0_APBmslave0_PADDR[0]), .Y(\sersta_m[4] ));
    SLE \sercon[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[0]_net_1 ));
    SLE \fsmsync[1]  (.D(N_955_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[1]_net_1 ));
    SLE \fsmmod[0]  (.D(\fsmmod_ns[0] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[0]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \SDAO_int_write_proc.un1_sersta65_1_0  
        (.A(\fsmsta[0]_net_1 ), .B(\fsmsta[1]_net_1 ), .C(N_1235), .D(
        sersta75), .Y(un1_sersta65_1_0));
    SLE \fsmmod[6]  (.D(N_1016_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[6]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \SDAI_ff_reg_proc.SDAI_ff_reg_3[1]  (.A(
        \sercon[6]_net_1 ), .B(\SDAI_ff_reg[0]_net_1 ), .Y(
        \SDAI_ff_reg_3[1] ));
    CFG4 #( .INIT(16'h0020) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_a4_1  (.A(
        counter_PRESETN_1_net_1), .B(fsmsta13), .C(adrcomp_net_1), .D(
        fsmsta33), .Y(N_1311));
    CFG4 #( .INIT(16'hDF00) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_a0_0  (.A(
        un1_framesync24_1_0), .B(sersta64), .C(adrcompen_net_1), .D(
        fsmsta_9_2_342_i_a4_0), .Y(fsmsta_9_2_342_i_a2_0));
    CFG3 #( .INIT(8'h51) )  fsmsta_nxt_1_sqmuxa_4_0 (.A(
        \fsmsta[0]_net_1 ), .B(\COREI2C_0_0_SDAO[0] ), .C(SDAInt_net_1)
        , .Y(fsmsta_nxt_1_sqmuxa_4_0_net_1));
    SLE \sercon[4]  (.D(\sercon_9[4] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sercon[4]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  \sersta_write_proc.sersta85  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(sersta85_1), .D(
        \fsmsta[1]_net_1 ), .Y(sersta85));
    CFG4 #( .INIT(16'h0040) )  \PRDATA_0_iv_RNO_0[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[1]), .B(COREI2C_0_0_INT[0]), .C(
        un1_PRDATA_1), .D(CoreAPB3_0_APBmslave0_PADDR[0]), .Y(
        \sercon_m[3] ));
    CFG3 #( .INIT(8'h31) )  \fsmsta_nxt_3_0_d_am[1]  (.A(N_7), .B(
        fsmsta_nxt93), .C(\fsmsta[1]_net_1 ), .Y(
        \fsmsta_nxt_3_0_d_am[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \sercon_write_proc.fsmmod_nxt_0_sqmuxa  (
        .A(\fsmmod[4]_net_1 ), .B(SCLInt_net_1), .C(PCLKint_p1_net_1), 
        .Y(fsmmod_nxt_0_sqmuxa));
    SLE SCLO_int (.D(SCLO_int5_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \COREI2C_0_0_SCLO[0] ));
    SLE \fsmmod[2]  (.D(N_1010_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[2]_net_1 ));
    CFG4 #( .INIT(16'h00E2) )  un1_fsmsta_nxt_1_sqmuxa_1_1 (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        fsmsta_nxt_1_sqmuxa_4_0_net_1), .D(\fsmsta[1]_net_1 ), .Y(
        un1_fsmsta_nxt_1_sqmuxa_1_1_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \un1_fsmsta_nxt_0_1_iv[1]  (.A(sersta65)
        , .B(sersta69), .C(\fsmsta_nxt_4_i_m[3] ), .D(
        \un1_fsmsta_nxt_0_1_iv_1[1]_net_1 ), .Y(\un1_fsmsta_nxt[1] ));
    SLE \sersta[3]  (.D(\sersta_3[3] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[3]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  \SDAO_int_write_proc.sersta72  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(sersta80_1), .D(
        \fsmsta[0]_net_1 ), .Y(sersta72));
    SLE \fsmsync[6]  (.D(N_965_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[6]_net_1 ));
    SLE \SDAI_ff_reg[2]  (.D(\SDAI_ff_reg_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[2]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  \sersta_write_proc.sersta66  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .D(\fsmsta[2]_net_1 ), .Y(sersta66));
    CFG4 #( .INIT(16'h7F40) )  
        \NoName_cnst_2_4_3__NoName_cnst_2_1_0_.m10  (.A(ack_net_1), .B(
        adrcompen_net_1), .C(un1_framesync24_1_0), .D(
        \fsmsta[3]_net_1 ), .Y(\NoName_cnst_2[3] ));
    SLE \fsmsync[0]  (.D(\fsmsync_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[0]_net_1 ));
    CFG4 #( .INIT(16'h5554) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_m4_s  (.A(un1_framesync24_0)
        , .B(un1_sersta84_2_0), .C(N_756), .D(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .Y(fsmsta_9_0_372_i_m4_s));
    SLE \PCLK_count1[0]  (.D(\PCLK_count1_4[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[0]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  \SDAO_int_write_proc.sersta61  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(N_1020_1), .Y(sersta61));
    CFG4 #( .INIT(16'h15D5) )  
        \NoName_cnst_2_4_3__NoName_cnst_2_1_0_.m4  (.A(N_4), .B(
        un1_framesync24_1_0), .C(adrcompen_net_1), .D(ack_net_1), .Y(
        N_5));
    CFG4 #( .INIT(16'hFBFA) )  \un1_fsmsta_nxt_0_0_iv[0]  (.A(sersta83)
        , .B(SDAInt_net_1), .C(\fsmsta_nxt_4_i_m[0] ), .D(
        un1_sersta60_net_1), .Y(\un1_fsmsta_nxt_0_0_iv[0]_net_1 ));
    CFG4 #( .INIT(16'hC8C0) )  \fsmsync_ns_0_a3_3[0]  (.A(
        \fsmmod[1]_net_1 ), .B(\fsmsync_ns_0_a3_3_0[0]_net_1 ), .C(
        \fsmmod[3]_net_1 ), .D(\fsmmod[2]_net_1 ), .Y(N_999));
    SLE \fsmsta[0]  (.D(\fsmsta_9[0] ), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\fsmsta[0]_net_1 ));
    SLE \serdat[3]  (.D(\serdat_19[3] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[3]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \fsmmod_ns_i_a4_1[2]  (.A(
        COREI2C_0_0_INT[0]), .B(\sercon[5]_net_1 ), .C(N_1059), .D(
        \fsmmod_ns_i_a4_0[2] ), .Y(\fsmmod_ns_i_a4_1[2]_net_1 ));
    CFG3 #( .INIT(8'h32) )  \fsmsta_sync_proc.fsmsta_9_bm[4]  (.A(
        ack_net_1), .B(\fsmsta_cnst_i_0[4]_net_1 ), .C(un1_fsmdet_0), 
        .Y(\fsmsta_9_bm[4] ));
    SLE nedetect (.D(nedetect_0_sqmuxa_net_1), .CLK(GL0_INST), .EN(
        SCLInt6), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        nedetect_net_1));
    CFG4 #( .INIT(16'hEEE2) )  \un1_SDAInt[2]  (.A(\fsmsta[2]_net_1 ), 
        .B(framesync24), .C(\sercon[2]_net_1 ), .D(SDAInt_net_1), .Y(
        N_1151));
    CFG4 #( .INIT(16'h3022) )  \serdat_write_proc.bsd7_tmp_7_ns  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .B(\fsmdet[3]_net_1 ), .C(
        bsd7_tmp_7_am), .D(bsd7_tmp_7_ns_1), .Y(bsd7_tmp_7));
    CFG4 #( .INIT(16'hFFEC) )  adrcompen_2_sqmuxa_i (.A(framesync24), 
        .B(adrcomp12), .C(nedetect_net_1), .D(\fsmdet[3]_net_1 ), .Y(
        adrcompen_2_sqmuxa_i_0));
    CFG2 #( .INIT(4'h4) )  \fsmmod_ns_0_a4_0_2[1]  (.A(fsmmod5), .B(
        \fsmmod[0]_net_1 ), .Y(N_1048_2));
    CFG4 #( .INIT(16'h1000) )  serdat_2_sqmuxa_1_0 (.A(
        COREI2C_0_0_INT[0]), .B(\fsmdet[3]_net_1 ), .C(un1_sersta58), 
        .D(\sercon[6]_net_1 ), .Y(serdat_2_sqmuxa_1_0_net_1));
    CFG4 #( .INIT(16'hF022) )  \sercon_write_proc.sercon_9[4]  (.A(
        \sercon_8_1[4] ), .B(un1_fsmdet_2_0), .C(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .D(sercon18), .Y(
        \sercon_9[4] ));
    CFG1 #( .INIT(2'h1) )  SCLO_int_RNI12J6 (.A(\COREI2C_0_0_SCLO[0] ), 
        .Y(COREI2C_0_0_SCLO_i[0]));
    CFG4 #( .INIT(16'hCCC6) )  
        \framesync_write_proc.framesync_6_enl_bm[0]  (.A(
        nedetect_net_1), .B(\framesync[0]_net_1 ), .C(framesync24), .D(
        un1_framesync_2), .Y(\framesync_6_enl_bm[0] ));
    CFG4 #( .INIT(16'h3ACA) )  
        \framesync_write_proc.framesync_6_enl[1]  (.A(
        \fsmdet[3]_net_1 ), .B(\framesync[1]_net_1 ), .C(
        framesync_6_e2), .D(CO0), .Y(\framesync_6[1] ));
    CFG4 #( .INIT(16'hCF9F) )  \sersta_write_proc.sersta_3[3]  (.A(
        sersta84_2), .B(\sersta_3_1[3] ), .C(COREI2C_0_0_INT[0]), .D(
        \fsmsta[3]_net_1 ), .Y(\sersta_3[3] ));
    CFG2 #( .INIT(4'hE) )  \fsmsync_ns_i_o3[3]  (.A(N_994), .B(
        COREI2C_0_0_INT[0]), .Y(N_973));
    CFG2 #( .INIT(4'h8) )  \SDAO_int_write_proc.sersta70_1  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(sersta85_1));
    CFG2 #( .INIT(4'hD) )  starto_en_1_sqmuxa_i (.A(starto_en8), .B(
        PCLKint_p1_net_1), .Y(starto_en_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'h0010) )  \SDAO_int_write_proc.sersta70  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(sersta85_1), .D(
        \fsmsta[1]_net_1 ), .Y(sersta70));
    CFG4 #( .INIT(16'hC888) )  un1_sersta84_2_1_0 (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .D(\fsmsta[1]_net_1 ), .Y(
        un1_sersta84_2_1_0_net_1));
    CFG3 #( .INIT(8'hE4) )  
        \framesync_write_proc.framesync_6_enl_ns[0]  (.A(
        framesync_6_e2), .B(\framesync_6_enl_am[0] ), .C(
        \framesync_6_enl_bm[0] ), .Y(\framesync_6[0] ));
    CFG3 #( .INIT(8'hFE) )  un1_sersta71 (.A(sersta71), .B(sersta75), 
        .C(sersta72), .Y(un1_sersta71_net_1));
    CFG3 #( .INIT(8'hD0) )  SDAO_int_1_sqmuxa_1 (.A(\fsmmod[0]_net_1 ), 
        .B(adrcomp_net_1), .C(N_1290_2), .Y(SDAO_int_1_sqmuxa_1_net_1));
    SLE \fsmsta[1]  (.D(N_1328_i_0), .CLK(GL0_INST), .EN(
        un1_ens1_pre_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\fsmsta[1]_net_1 ));
    CFG4 #( .INIT(16'hF2F0) )  \serdat_write_proc.bsd7_tmp_7_am  (.A(
        un1_sersta58), .B(serdat4), .C(bsd7_tmp_net_1), .D(
        bsd7_tmp_7_sn_m6_1_0), .Y(bsd7_tmp_7_am));
    CFG3 #( .INIT(8'h08) )  SDAO_int_1_sqmuxa_2 (.A(\sercon[6]_net_1 ), 
        .B(N_1290_1), .C(\fsmmod[3]_net_1 ), .Y(
        SDAO_int_1_sqmuxa_2_net_1));
    CFG3 #( .INIT(8'h04) )  \fsmmod_ns_0_a4[1]  (.A(fsmmod5), .B(
        \fsmmod[1]_net_1 ), .C(nedetect_net_1), .Y(N_1040));
    CFG4 #( .INIT(16'h0010) )  un1_fsmdet_1_2 (.A(\fsmdet[5]_net_1 ), 
        .B(PCLK_count2_ov_net_1), .C(N_827), .D(\fsmdet[3]_net_1 ), .Y(
        un1_fsmdet_1_2_net_1));
    CFG3 #( .INIT(8'h06) )  un1_sersta60 (.A(\fsmsta[2]_net_1 ), .B(
        \fsmsta[1]_net_1 ), .C(N_1020_1), .Y(un1_sersta60_net_1));
    CFG2 #( .INIT(4'h1) )  \serdat_write_proc.bsd7_10_iv_i_1_RNO  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .B(COREI2C_0_0_INT[0]), .Y(
        \PWDATA_i_m_0[7] ));
    CFG4 #( .INIT(16'h1000) )  \SDAO_int_write_proc.sersta69  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(N_1236_2), .Y(sersta69));
    SLE \SDAI_ff_reg[3]  (.D(\SDAI_ff_reg_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[3]_net_1 ));
    CFG4 #( .INIT(16'h48C0) )  \PCLK_counter1_proc.PCLK_count1_4[3]  (
        .A(CO1), .B(PCLK_count1_0_sqmuxa_net_1), .C(
        \PCLK_count1[3]_net_1 ), .D(\PCLK_count1[2]_net_1 ), .Y(
        \PCLK_count1_4[3] ));
    CFG4 #( .INIT(16'hFF15) )  
        \framesync_write_proc.framesync_6_enl_am[0]  (.A(framesync10), 
        .B(framesync14), .C(un1_framesync_2), .D(framesync_6_sm0), .Y(
        \framesync_6_enl_am[0] ));
    SLE \framesync[0]  (.D(\framesync_6[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \framesync[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \SDAO_int_write_proc.sersta64_1  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[2]_net_1 ), .Y(sersta80_1));
    SLE bsd7_tmp (.D(bsd7_tmp_7), .CLK(GL0_INST), .EN(
        \sercon[6]_net_1 ), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(bsd7_tmp_net_1));
    SLE \fsmdet[3]  (.D(N_875_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[3]_net_1 ));
    CFG3 #( .INIT(8'h01) )  un1_counter_PRESETN_i_a2 (.A(
        \fsmsync[1]_net_1 ), .B(\fsmsync[5]_net_1 ), .C(
        \fsmsync[4]_net_1 ), .Y(N_827));
    SLE PCLKint_ff (.D(PCLKint_ff_3), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PCLKint_ff_net_1));
    SLE \serdat[6]  (.D(\serdat_19[6] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \fsmdet_RNO[0]  (.A(SCLInt_net_1), .Y(
        SCLInt_i_0));
    CFG4 #( .INIT(16'h0111) )  \fsmmod_RNO[2]  (.A(
        \fsmmod_ns_i_0_0[2]_net_1 ), .B(fsmmod5), .C(
        \fsmmod_ns_i_a4_1[2]_net_1 ), .D(\fsmmod_ns_i_a4_2[2]_net_1 ), 
        .Y(N_1010_i_0));
    CFG3 #( .INIT(8'hF1) )  \un1_fsmsta_nxt_1[3]  (.A(
        \un1_fsmsta_nxt_0_1_iv[3]_net_1 ), .B(un1_sersta84_1_1_0_net_1)
        , .C(un1_sersta84_1_2_net_1), .Y(\un1_fsmsta_nxt_1[3]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \fsmsta_sync_proc.un1_fsmdet  (.A(
        counter_PRESETN_1_net_1), .B(fsmsta33), .Y(un1_fsmdet_0));
    CFG4 #( .INIT(16'h0200) )  \SDAO_int_write_proc.sersta78_3  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(\fsmsta[2]_net_1 ), .Y(sersta78_3));
    CFG2 #( .INIT(4'h8) )  \fsmsync_sync_proc.un1_sersta69_1_a5_2  (.A(
        N_1237_2), .B(N_1237_1), .Y(N_1237));
    CFG4 #( .INIT(16'h000B) )  \fsmmod_RNO[6]  (.A(\fsmmod[3]_net_1 ), 
        .B(nedetect_net_1), .C(N_1049), .D(fsmmod5), .Y(N_1016_i_0));
    CFG3 #( .INIT(8'h02) )  un1_sersta84_2_1_a6_1 (.A(framesync24), .B(
        sersta80_1), .C(N_1020_1), .Y(N_1225));
    CFG4 #( .INIT(16'h1373) )  \sersta_write_proc.sersta_2_4_0_.m21  (
        .A(\fsmsta[2]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(\fsmsta[0]_net_1 ), .Y(N_22));
    CFG3 #( .INIT(8'h40) )  \SDAO_int_write_proc.sersta73_0  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[3]_net_1 ), .Y(N_1235));
    SLE bsd7 (.D(bsd7_10_iv_i_0), .CLK(GL0_INST), .EN(
        \sercon[6]_net_1 ), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(bsd7_net_1));
    SLE PCLKint (.D(PCLKint_4), .CLK(GL0_INST), .EN(un1_fsmdet_1_i_0), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PCLKint_net_1));
    SLE \PCLK_count1[1]  (.D(\PCLK_count1_4[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[1]_net_1 ));
    SLE \serdat[5]  (.D(\serdat_19[5] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[5]_net_1 ));
    CFG4 #( .INIT(16'hECCC) )  \fsmsync_ns_0[0]  (.A(N_972), .B(
        \fsmsync_ns_0_1[0]_net_1 ), .C(\fsmsync[0]_net_1 ), .D(
        SCLInt_net_1), .Y(\fsmsync_ns[0] ));
    CFG4 #( .INIT(16'h0D00) )  fsmsta_3_sqmuxa_0 (.A(un1_framesync_4), 
        .B(COREI2C_0_0_INT[0]), .C(un1_fsmsta33), .D(
        counter_PRESETN_1_net_1), .Y(fsmsta_3_sqmuxa_0_net_1));
    CFG4 #( .INIT(16'hF3F1) )  \fsmmod_ns_i_0_0[2]  (.A(nedetect_net_1)
        , .B(\fsmmod[2]_net_1 ), .C(N_1052), .D(N_1059), .Y(
        \fsmmod_ns_i_0_0[2]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_0_iv[5]  (.A(\serdat[5]_net_1 ), 
        .B(\sersta_m[2] ), .C(\sercon_m[5] ), .D(un4_PRDATA), .Y(
        \PRDATAi[0]_4 ));
    CFG3 #( .INIT(8'h80) )  \SDAO_int_write_proc.sersta65  (.A(
        \fsmsta[1]_net_1 ), .B(sersta65_1), .C(\fsmsta[0]_net_1 ), .Y(
        sersta65));
    CFG2 #( .INIT(4'h1) )  SDAO_int_1_sqmuxa_5 (.A(\fsmmod[4]_net_1 ), 
        .B(\fsmmod[6]_net_1 ), .Y(N_1290_2));
    CFG3 #( .INIT(8'h01) )  \PRDATA_0_iv_RNO_1[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[0]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        \PRDATA_0_iv_RNO_1[7]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \adrcomp_write_proc.un1_sercon_1_4  (.A(
        \serdat[5]_net_1 ), .B(serdat_4), .C(\serdat[3]_net_1 ), .D(
        nedetect_net_1), .Y(un1_sercon_1_4));
    CFG2 #( .INIT(4'hE) )  \framesync_write_proc.framesync_6s2  (.A(
        counter_PRESETN_1_net_1), .B(bsd7_tmp_i_m_1), .Y(
        framesync_6_sm0));
    CFG2 #( .INIT(4'h7) )  \sersta_write_proc.sersta_3[2]  (.A(
        N_26_mux), .B(COREI2C_0_0_INT[0]), .Y(\sersta_3[2] ));
    CFG4 #( .INIT(16'h0405) )  \fsmsync_RNO[4]  (.A(SCLInt_net_1), .B(
        \fsmsync[4]_net_1 ), .C(N_985), .D(N_980), .Y(N_961_i_0));
    CFG4 #( .INIT(16'h0100) )  \adrcomp_write_proc.fsmsta19  (.A(
        \serdat[6]_net_1 ), .B(\serdat[5]_net_1 ), .C(
        \serdat[1]_net_1 ), .D(fsmsta19_2_0), .Y(fsmsta19));
    SLE \SDAI_ff_reg[0]  (.D(\SDAI_ff_reg_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \fsmsync_RNO[5]  (.A(COREI2C_0_0_INT[0]), 
        .B(N_994), .C(N_985), .Y(N_963_i_0));
    CFG4 #( .INIT(16'hAAA3) )  \un1_fsmsta_nxt_1[0]  (.A(
        \fsmsta[0]_net_1 ), .B(\un1_fsmsta_nxt_0_0_iv[0]_net_1 ), .C(
        un1_sersta84_1_1_0_net_1), .D(un1_sersta84_1_2_net_1), .Y(
        \un1_fsmsta_nxt_1[0]_net_1 ));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[6]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .B(\serdat[5]_net_1 ), .C(
        un1_PSEL), .D(un4_PRDATA), .Y(\serdat_19[6] ));
    CFG4 #( .INIT(16'hFFFE) )  \fsmmod_ns_i_o4_1[2]  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(\fsmsta[2]_net_1 ), .Y(N_1020));
    SLE adrcomp (.D(un1_adrcomp14_1_net_1), .CLK(GL0_INST), .EN(
        adrcomp_2_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(adrcomp_net_1));
    CFG3 #( .INIT(8'h80) )  \adrcomp_write_proc.sersta81  (.A(
        \fsmsta[1]_net_1 ), .B(sersta81_0), .C(\fsmsta[0]_net_1 ), .Y(
        sersta81));
    CFG4 #( .INIT(16'h4000) )  \adrcomp_write_proc.sersta77_3  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .D(\fsmsta[1]_net_1 ), .Y(sersta77_3));
    CFG2 #( .INIT(4'hE) )  \PCLKint_write_proc.PCLKint_ff_3  (.A(
        counter_PRESETN), .B(PCLKint_net_1), .Y(PCLKint_ff_3));
    CFG2 #( .INIT(4'hE) )  \fsmsta_cnst_0_o4[2]  (.A(fsmsta19), .B(
        ack_net_1), .Y(N_1072));
    CFG4 #( .INIT(16'h23AF) )  \serdat_write_proc.bsd7_10_iv_i_1  (.A(
        bsd7_net_1), .B(\PWDATA_i_m_0[7] ), .C(
        \un1_bsd7_1_sqmuxa[0]_net_1 ), .D(serdat4), .Y(bsd7_10_iv_i_1));
    SLE adrcompen (.D(un1_adrcomp14_net_1), .CLK(GL0_INST), .EN(
        adrcompen_2_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(adrcompen_net_1));
    CFG4 #( .INIT(16'hF0F1) )  \fsmsync_ns_i_0[3]  (.A(
        \fsmsync[2]_net_1 ), .B(\fsmsync[5]_net_1 ), .C(N_985), .D(
        N_974), .Y(\fsmsync_ns_i_0[3]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  \fsmsta_sync_proc.un1_framesync24  (.A(
        pedetect_net_1), .B(adrcompen_net_1), .C(un1_framesync24_1_0), 
        .D(sersta64), .Y(un1_framesync24_0));
    CFG3 #( .INIT(8'hD8) )  \fsmsta_nxt_3[0]  (.A(un1_sersta84_2_0), 
        .B(\un1_fsmsta_nxt_1[0]_net_1 ), .C(N_1126), .Y(
        \fsmsta_nxt_3[0]_net_1 ));
    SLE \SDAI_ff_reg[1]  (.D(\SDAI_ff_reg_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SDAI_ff_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[1]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .B(serdat_0), .C(un1_PSEL), 
        .D(un4_PRDATA), .Y(\serdat_19[1] ));
    CFG2 #( .INIT(4'h8) )  \adrcomp_write_proc.sersta83_0  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(sersta84_2));
    CFG3 #( .INIT(8'h80) )  \sercon_write_proc.un1_PRDATA_1_RNIVTQD  (
        .A(un1_PRDATA_1), .B(\sercon[4]_net_1 ), .C(un14_PRDATA_2), .Y(
        sercon_m_4));
    CFG4 #( .INIT(16'h2000) )  PCLK_count2_ov_0_sqmuxa (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN), .C(
        \PCLK_count2[1]_net_1 ), .D(\PCLK_count2[0]_net_1 ), .Y(
        PCLK_count2_ov_0_sqmuxa_net_1));
    SLE \fsmdet[6]  (.D(N_881_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[6]_net_1 ));
    CFG4 #( .INIT(16'hFFF2) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_1_1  
        (.A(un1_fsmmod_1), .B(fsmsta33), .C(fsmsta_9_2_342_i_a3), .D(
        N_1311), .Y(fsmsta_9_2_342_i_1_1));
    CFG3 #( .INIT(8'hF7) )  \fsmmod_ns_0_o4[0]  (.A(starto_en_net_1), 
        .B(PCLKint_p1_net_1), .C(N_1029), .Y(N_1031));
    CFG3 #( .INIT(8'h7F) )  \fsmsync_ns_i_o3[4]  (.A(
        \indelay[1]_net_1 ), .B(\indelay[2]_net_1 ), .C(
        \fsmsync[3]_net_1 ), .Y(N_980));
    CFG4 #( .INIT(16'hAAEA) )  \fsmmod_ns_0[1]  (.A(N_1040), .B(
        N_1048_2), .C(SDAInt_net_1), .D(N_1031), .Y(\fsmmod_ns[1] ));
    CFG3 #( .INIT(8'h08) )  \adrcomp_write_proc.sersta81_0  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[3]_net_1 ), .Y(sersta81_0));
    CFG4 #( .INIT(16'h8000) )  ack_bit_1_sqmuxa (.A(serdat48), .B(
        sercon18), .C(COREI2C_0_0_INT[0]), .D(\sercon[6]_net_1 ), .Y(
        ack_bit_1_sqmuxa_net_1));
    CFG2 #( .INIT(4'h1) )  pedetect_0_sqmuxa (.A(SCLInt6), .B(
        SCLInt_net_1), .Y(pedetect_0_sqmuxa_net_1));
    CFG2 #( .INIT(4'h1) )  mst_0_a2 (.A(\fsmmod[5]_net_1 ), .B(
        \fsmmod[0]_net_1 ), .Y(mst));
    CFG4 #( .INIT(16'hFFFE) )  \un1_fsmsta_nxt_0_1_iv[3]  (.A(sersta75)
        , .B(\fsmsta_nxt_4_i_m[3] ), .C(sersta65), .D(
        un1_sersta60_net_1), .Y(\un1_fsmsta_nxt_0_1_iv[3]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \SDAO_int_write_proc.un1_sersta65_1  (.A(
        un1_sersta65_1_1_0), .B(un1_sersta65_1_0), .C(un1_sersta65_1_1)
        , .Y(un1_sersta65_1));
    CFG4 #( .INIT(16'h0004) )  \SDAO_int_write_proc.framesync24  (.A(
        \framesync[2]_net_1 ), .B(\framesync[3]_net_1 ), .C(
        \framesync[1]_net_1 ), .D(\framesync[0]_net_1 ), .Y(
        framesync24));
    SLE \sersta[4]  (.D(\sersta_3[4] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[4]_net_1 ));
    SLE SCLInt (.D(\SCLI_ff_reg[3]_net_1 ), .CLK(GL0_INST), .EN(
        un1_SCLInt5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        SCLInt_net_1));
    CFG4 #( .INIT(16'h0B0F) )  
        \fsmsta_sync_proc.fsmsta_9_2_342_i_a4_0_0  (.A(PCLKint_net_1), 
        .B(PCLKint_ff_net_1), .C(counter_PRESETN_1_net_1), .D(
        \fsmmod[4]_net_1 ), .Y(fsmsta_9_2_342_i_a4_0));
    CFG3 #( .INIT(8'hE2) )  \fsmsta_nxt_3_0_d_ns[1]  (.A(
        \fsmsta_nxt_3_0_d_am[1]_net_1 ), .B(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .C(
        \fsmsta_nxt_3_0_d_bm[1]_net_1 ), .Y(
        \fsmsta_nxt_3_0_d_ns[1]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  un1_serdat_2_sqmuxa (.A(
        serdat_2_sqmuxa_1_0_net_1), .B(pedetect_net_1), .C(serdat4), 
        .D(un1_serdat_2_sqmuxa_1_1_net_1), .Y(
        un1_serdat_2_sqmuxa_net_1));
    CFG4 #( .INIT(16'h8DA5) )  \un1_fsmsta_nxt_2_ns[4]  (.A(
        un1_fsmsta_nxt_2_sn_N_3), .B(\COREI2C_0_0_SDAO[0] ), .C(
        \un1_fsmsta_nxt_2_ns_1[4]_net_1 ), .D(un1_framesync24_1_net_1), 
        .Y(N_1124));
    CFG2 #( .INIT(4'h7) )  \sersta_write_proc.sersta_3[1]  (.A(
        N_25_mux), .B(COREI2C_0_0_INT[0]), .Y(\sersta_3[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \SDAO_int_write_proc.un1_sersta65_1_1_0  (.A(sersta71), .B(
        sersta67), .C(sersta65), .D(sersta72), .Y(un1_sersta65_1_1_0));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_RNO_0[7]  (.A(
        \PRDATA_0_iv_RNO_1[7]_net_1 ), .B(\sercon[7]_net_1 ), .C(
        un14_PRDATA_net_1), .D(un9_PRDATA_2_0), .Y(\PRDATA_0_iv_0[7] ));
    SLE PCLK_count2_ov (.D(PCLK_count2_ov_0_sqmuxa_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PCLK_count2_ov_net_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA_0_iv_RNO_0[5]  (.A(un1_PRDATA_1), 
        .B(\sercon[5]_net_1 ), .C(un14_PRDATA_2), .Y(\sercon_m[5] ));
    CFG2 #( .INIT(4'h4) )  un1_adrcomp14 (.A(adrcomp12), .B(
        \fsmdet[3]_net_1 ), .Y(un1_adrcomp14_net_1));
    CFG4 #( .INIT(16'h0080) )  \PRDATA_0_iv_RNO[5]  (.A(
        un9_PRDATA_1_net_1), .B(un9_PRDATA_2_0), .C(\sersta[2]_net_1 ), 
        .D(CoreAPB3_0_APBmslave0_PADDR[0]), .Y(\sersta_m[2] ));
    CFG2 #( .INIT(4'hE) )  \busfree_write_proc.un1_fsmdet_2  (.A(
        adrcomp12), .B(\fsmdet[5]_net_1 ), .Y(un1_fsmdet_2_0));
    CFG2 #( .INIT(4'h8) )  \un1_framesync_1_1.CO1  (.A(CO0), .B(
        \framesync[1]_net_1 ), .Y(CO1_0));
    CFG4 #( .INIT(16'h0103) )  \fsmsync_RNO[2]  (.A(\fsmsync[0]_net_1 )
        , .B(N_989), .C(N_985), .D(N_983), .Y(N_957_i_0));
    SLE \sercon[3]  (.D(\sercon_9[3] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        COREI2C_0_0_INT[0]));
    CFG3 #( .INIT(8'hF1) )  \sercon_write_proc.un1_adrcomp  (.A(
        \fsmmod[5]_net_1 ), .B(\fsmmod[0]_net_1 ), .C(adrcomp_net_1), 
        .Y(un1_adrcomp));
    CFG3 #( .INIT(8'h01) )  \sercon_write_proc.un1_PRDATA_1_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(un1_PRDATA_1));
    SLE \fsmmod[5]  (.D(\fsmmod_ns[5] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \adrcomp_write_proc.sersta77  (.A(
        sersta77_3), .B(\fsmsta[2]_net_1 ), .Y(sersta77));
    CFG4 #( .INIT(16'h0001) )  \adrcomp_write_proc.fsmsta19_2_0  (.A(
        serdat_4), .B(\serdat[3]_net_1 ), .C(\serdat[2]_net_1 ), .D(
        serdat_0), .Y(fsmsta19_2_0));
    CFG3 #( .INIT(8'h74) )  SDAO_int_1_sqmuxa_4_0 (.A(nedetect_net_1), 
        .B(un1_framesync_1), .C(framesync24), .Y(
        SDAO_int_1_sqmuxa_4_net_1));
    CFG3 #( .INIT(8'h40) )  un1_serdat_2_sqmuxa_1 (.A(serdat4), .B(
        pedetect_net_1), .C(un1_serdat_2_sqmuxa_1_tz_net_1), .Y(
        un1_serdat_2_sqmuxa_1_net_1));
    CFG2 #( .INIT(4'h1) )  \PCLK_counter1_proc.PCLK_count1_ov_3  (.A(
        counter_PRESETN), .B(PCLK_count17), .Y(PCLK_count1_ov_3));
    CFG3 #( .INIT(8'hEF) )  \fsmmod_ns_0_o3[3]  (.A(\sercon[4]_net_1 ), 
        .B(COREI2C_0_0_INT[0]), .C(\sercon[5]_net_1 ), .Y(N_1029));
    CFG4 #( .INIT(16'h00C8) )  un1_sersta84_2_1_a6_0 (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(sersta80_1), .D(
        framesync24), .Y(N_1224));
    CFG4 #( .INIT(16'h4044) )  un1_fsmsta_nxt_1_sqmuxa_1 (.A(N_1020_1), 
        .B(un1_fsmsta_nxt_1_sqmuxa_1_1_net_1), .C(\fsmsta[2]_net_1 ), 
        .D(fsmsta_nxt19), .Y(un1_fsmsta_nxt_1_sqmuxa_1_net_1));
    CFG2 #( .INIT(4'h8) )  un1_framesync24_1 (.A(un1_sersta69_net_1), 
        .B(framesync24), .Y(un1_framesync24_1_net_1));
    CFG3 #( .INIT(8'h10) )  un18_counter_PRESETN (.A(SCLInt_net_1), .B(
        \fsmmod[5]_net_1 ), .C(busfree_net_1), .Y(
        un18_counter_PRESETN_net_1));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[7]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .B(\serdat[6]_net_1 ), .C(
        un1_PSEL), .D(un4_PRDATA), .Y(\serdat_19[7] ));
    SLE \fsmdet[5]  (.D(N_879_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmdet[5]_net_1 ));
    SLE \fsmmod[1]  (.D(\fsmmod_ns[1] ), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmmod[1]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  \sersta_RNIIFT31[3]  (.A(
        un9_PRDATA_1_net_1), .B(un9_PRDATA_2_0), .C(\sersta[3]_net_1 ), 
        .D(CoreAPB3_0_APBmslave0_PADDR[0]), .Y(sersta_m_3));
    CFG4 #( .INIT(16'hAE00) )  \fsmdet_RNO[4]  (.A(\fsmdet[3]_net_1 ), 
        .B(\fsmdet[4]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_877_i_0));
    CFG4 #( .INIT(16'hE000) )  \fsmdet_RNO[1]  (.A(\fsmdet[0]_net_1 ), 
        .B(\fsmdet[1]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_871_i_0));
    CFG4 #( .INIT(16'h4F7F) )  \sersta_write_proc.sersta_3[0]  (.A(
        N_4_0), .B(sersta84_2), .C(COREI2C_0_0_INT[0]), .D(
        \fsmsta[0]_net_1 ), .Y(\sersta_3[0] ));
    CFG4 #( .INIT(16'hFFFE) )  un1_sersta84_1_2 (.A(sersta85), .B(
        sersta66), .C(sersta82), .D(sersta84), .Y(
        un1_sersta84_1_2_net_1));
    SLE \fsmsync[4]  (.D(N_961_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[4]_net_1 ));
    CFG3 #( .INIT(8'h70) )  
        \fsmsta_sync_proc.fsmsta_9_0_372_i_m4_s_RNO  (.A(framesync24), 
        .B(un1_sersta69_net_1), .C(un1_fsmsta_nxt_2_sn_N_3), .Y(N_756));
    CFG3 #( .INIT(8'hFE) )  un1_sersta84_1_1_0 (.A(sersta76), .B(
        sersta77_3), .C(sersta74), .Y(un1_sersta84_1_1_0_net_1));
    CFG3 #( .INIT(8'hE0) )  \fsmsta_cnst_i_0[4]  (.A(\fsmmod[6]_net_1 )
        , .B(\fsmmod[1]_net_1 ), .C(\fsmdet[3]_net_1 ), .Y(
        \fsmsta_cnst_i_0[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \sercon_RNIRPQD[0]  (.A(un1_PRDATA_1), .B(
        \sercon[0]_net_1 ), .C(un14_PRDATA_2), .Y(sercon_m_0));
    CFG2 #( .INIT(4'hD) )  sclscl_1_sqmuxa_i (.A(\fsmmod[5]_net_1 ), 
        .B(pedetect_net_1), .Y(sclscl_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'hFEFA) )  \PRDATA_0_iv[7]  (.A(\sersta_m[4] ), .B(
        \serdat[7]_net_1 ), .C(\PRDATA_0_iv_0[7] ), .D(un4_PRDATA), .Y(
        \PRDATAi[0]_6 ));
    CFG4 #( .INIT(16'h0054) )  \fsmsta_RNO[3]  (.A(
        fsmsta_9_2_342_i_1_1), .B(un1_sersta84_2_0), .C(N_1306_i_1), 
        .D(fsmsta_9_2_342_i_a2), .Y(N_1306_i_0));
    SLE \sercon[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[5]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  \adrcomp_write_proc.sersta82  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(N_1237_2), .D(
        \fsmsta[1]_net_1 ), .Y(sersta82));
    CFG2 #( .INIT(4'h2) )  SCLInt_RNIEO25 (.A(COREI2C_0_0_INT[0]), .B(
        SCLInt_net_1), .Y(bsd7_tmp_i_m_1));
    CFG4 #( .INIT(16'h008A) )  \fsmsync_ns_i_a3[3]  (.A(
        \sercon[4]_net_1 ), .B(un1_framesync_2), .C(\fsmsync[2]_net_1 )
        , .D(\fsmsync[3]_net_1 ), .Y(N_990));
    CFG3 #( .INIT(8'h08) )  \sercon_write_proc.sercon_8_1[4]  (.A(
        \sercon[4]_net_1 ), .B(\sercon[6]_net_1 ), .C(fsmsta33), .Y(
        \sercon_8_1[4] ));
    CFG3 #( .INIT(8'h7F) )  \serdat_write_proc.bsd7_tmp_7_ns_1  (.A(
        serdat4), .B(COREI2C_0_0_INT[0]), .C(un1_sersta58), .Y(
        bsd7_tmp_7_ns_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA_0_iv_RNO[2]  (.A(un1_PRDATA_1), .B(
        \sercon[2]_net_1 ), .C(un14_PRDATA_2), .Y(\sercon_m[2] ));
    CFG3 #( .INIT(8'h10) )  \PCLK_counter1_proc.PCLK_count1_4[0]  (.A(
        counter_PRESETN), .B(\PCLK_count1[0]_net_1 ), .C(PCLK_count17), 
        .Y(\PCLK_count1_4[0] ));
    CFG4 #( .INIT(16'h2220) )  serdat_0_sqmuxa (.A(COREI2C_0_0_INT[0]), 
        .B(\fsmdet[3]_net_1 ), .C(un1_sersta58_1), .D(
        un1_sersta60_1_net_1), .Y(serdat_0_sqmuxa_net_1));
    CFG3 #( .INIT(8'h62) )  \sersta_write_proc.sersta_2_4_0_.m3  (.A(
        \fsmsta[1]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[0]_net_1 ), .Y(N_4_0));
    CFG2 #( .INIT(4'h7) )  \SCLInt_write_proc.un1_SCLInt5  (.A(
        un1_SCLI_ff_reg), .B(SCLInt6), .Y(un1_SCLInt5));
    CFG4 #( .INIT(16'h000B) )  \fsmmod_RNO[4]  (.A(un1_framesync_2), 
        .B(\fsmmod[2]_net_1 ), .C(fsmmod5), .D(
        \fsmmod_ns_i_0[4]_net_1 ), .Y(N_1013_i_0));
    CFG4 #( .INIT(16'hFFFE) )  \SCLInt_write_proc.un1_SCLI_ff_reg  (.A(
        \SCLI_ff_reg[0]_net_1 ), .B(\SCLI_ff_reg[3]_net_1 ), .C(
        \SCLI_ff_reg[2]_net_1 ), .D(\SCLI_ff_reg[1]_net_1 ), .Y(
        un1_SCLI_ff_reg));
    SLE \SCLI_ff_reg[2]  (.D(\SCLI_ff_reg_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \SCLI_ff_reg[2]_net_1 ));
    CFG4 #( .INIT(16'hB0C0) )  \indelay_4[1]  (.A(\indelay[2]_net_1 ), 
        .B(\indelay[0]_net_1 ), .C(\fsmsync[3]_net_1 ), .D(
        \indelay[1]_net_1 ), .Y(\indelay_4[1]_net_1 ));
    CFG4 #( .INIT(16'h0031) )  \fsmsync_RNO[3]  (.A(N_973), .B(
        \fsmsync_ns_i_0[3]_net_1 ), .C(\fsmsync[3]_net_1 ), .D(N_990), 
        .Y(N_959_i_0));
    SLE \fsmsync[3]  (.D(N_959_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[3]_net_1 ));
    CFG4 #( .INIT(16'h3FAF) )  \sersta_write_proc.sersta_3[4]  (.A(
        \fsmsta[4]_net_1 ), .B(N_22), .C(COREI2C_0_0_INT[0]), .D(
        \fsmsta[3]_net_1 ), .Y(\sersta_3[4] ));
    CFG4 #( .INIT(16'h0103) )  \SDAO_int_write_proc.sersta67_RNI3QRD1  
        (.A(framesync24), .B(sersta65), .C(sersta67), .D(
        un1_sersta71_net_1), .Y(un1_fsmsta_nxt_2_sn_N_3));
    SLE \PCLK_count2[1]  (.D(\PCLK_count2_4[1]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\PCLK_count2[1]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  \serdat_write_proc.un4_PRDATA  (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(psh_enable_reg1_1_sqmuxa_0)
        , .C(CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(un4_PRDATA));
    CFG4 #( .INIT(16'h1230) )  \PCLK_count2_4[1]  (.A(
        PCLK_count1_ov_net_1), .B(counter_PRESETN), .C(
        \PCLK_count2[1]_net_1 ), .D(\PCLK_count2[0]_net_1 ), .Y(
        \PCLK_count2_4[1]_net_1 ));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[3]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .B(\serdat[2]_net_1 ), .C(
        un1_PSEL), .D(un4_PRDATA), .Y(\serdat_19[3] ));
    CFG4 #( .INIT(16'hA8A0) )  \sercon_write_proc.un1_fsmmod_2_2  (.A(
        un1_adrcomp), .B(un1_framesync24), .C(un1_sersta64_0), .D(
        counter_PRESETN_1_net_1), .Y(un1_fsmmod_2_2));
    CFG2 #( .INIT(4'h8) )  \fsmmod_ns_i_a4_2[2]  (.A(N_1020), .B(
        un1_framesync_2), .Y(\fsmmod_ns_i_a4_2[2]_net_1 ));
    CFG4 #( .INIT(16'h1A95) )  \sersta_write_proc.sersta_2_4_0_.m11  (
        .A(\fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(sersta84_2), 
        .D(\fsmsta[1]_net_1 ), .Y(N_25_mux));
    CFG4 #( .INIT(16'h0600) )  \PCLK_counter1_proc.PCLK_count1_4[2]  (
        .A(CO1), .B(\PCLK_count1[2]_net_1 ), .C(counter_PRESETN), .D(
        PCLK_count17), .Y(\PCLK_count1_4[2] ));
    CFG2 #( .INIT(4'h1) )  \fsmsync_ns_0_a3_3_0[0]  (.A(
        \fsmmod[5]_net_1 ), .B(\fsmmod[6]_net_1 ), .Y(
        \fsmsync_ns_0_a3_3_0[0]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \sercon_write_proc.un1_PRDATA_1  (.A(
        CoreAPB3_0_APBmslave0_PADDR[0]), .B(
        CoreAPB3_0_APBmslave0_PADDR[1]), .Y(un14_PRDATA_2));
    SLE busfree (.D(\fsmdet_i_0[3] ), .CLK(GL0_INST), .EN(un1_fsmdet), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(busfree_net_1));
    CFG3 #( .INIT(8'hD8) )  
        \framesync_write_proc.framesync_6_enl_ns[3]  (.A(
        framesync_6_e2), .B(\framesync_6_enl_bm[3] ), .C(
        \framesync_6_enl_am[3] ), .Y(\framesync_6[3] ));
    CFG3 #( .INIT(8'h20) )  \starto_en_write_proc.starto_en8  (.A(
        SCLInt_net_1), .B(\fsmmod[5]_net_1 ), .C(busfree_net_1), .Y(
        starto_en8));
    CFG2 #( .INIT(4'hD) )  \SMBint_filter_proc.SCLI_ff_reg_3[3]  (.A(
        \sercon[6]_net_1 ), .B(\SCLI_ff_reg[2]_net_1 ), .Y(
        \SCLI_ff_reg_3[3] ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_0_iv[2]  (.A(\serdat[2]_net_1 ), 
        .B(un14_PRDATA_net_1), .C(\sercon_m[2] ), .D(un4_PRDATA), .Y(
        \PRDATAi[0]_1 ));
    SLE \PCLK_count1[2]  (.D(\PCLK_count1_4[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \PCLK_count1[2]_net_1 ));
    CFG4 #( .INIT(16'hCCCD) )  \fsmsync_ns_i_1[6]  (.A(un1_framesync_2)
        , .B(\fsmsync_ns_i_0[6]_net_1 ), .C(\fsmsync[6]_net_1 ), .D(
        \fsmsync[5]_net_1 ), .Y(\fsmsync_ns_i_1[6]_net_1 ));
    SLE \sercon[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(sercon18), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sercon[6]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \SDAO_int_write_proc.sersta65_1  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[3]_net_1 ), .Y(sersta65_1));
    SLE SDAO_int (.D(N_1272), .CLK(GL0_INST), .EN(
        SDAO_int_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\COREI2C_0_0_SDAO[0] ));
    CFG4 #( .INIT(16'hFDDD) )  \fsmmod_sync_proc.fsmmod5  (.A(
        \sercon[6]_net_1 ), .B(\fsmdet[5]_net_1 ), .C(sersta64), .D(
        un1_sersta64_0), .Y(fsmmod5));
    CFG4 #( .INIT(16'hEAAA) )  \SDAO_int_write_proc.SDAO_int_6_0_312  
        (.A(SDAO_int_6_0_312_1), .B(N_1289), .C(N_1290_2), .D(N_1290_1)
        , .Y(N_1272));
    CFG3 #( .INIT(8'h07) )  \un1_fsmsta_nxt_2_am[3]  (.A(framesync24), 
        .B(un1_sersta71_net_1), .C(fsmsta_nxt19), .Y(
        \un1_fsmsta_nxt_2_am[3]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  \SDAO_int_write_proc.sersta71  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[3]_net_1 ), .C(un1_fsmsta), .D(
        \fsmsta[1]_net_1 ), .Y(sersta71));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[2]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .B(\serdat[1]_net_1 ), .C(
        un1_PSEL), .D(un4_PRDATA), .Y(\serdat_19[2] ));
    CFG4 #( .INIT(16'h2000) )  \adrcomp_write_proc.sersta76  (.A(
        \fsmsta[4]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(sersta74_2), .Y(sersta76));
    CFG3 #( .INIT(8'hB8) )  \fsmsta_nxt_3_RNO[0]  (.A(N_1149), .B(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .C(\un1_fsmsta_nxt_2[0] ), .Y(
        N_1126));
    CFG3 #( .INIT(8'h70) )  \un1_fsmsta_nxt_2_0[2]  (.A(framesync24), 
        .B(un1_sersta71_net_1), .C(fsmsta_nxt19), .Y(N_1110));
    CFG4 #( .INIT(16'h0020) )  \SDAO_int_write_proc.sersta64  (.A(
        \fsmsta[2]_net_1 ), .B(\fsmsta[0]_net_1 ), .C(
        \fsmsta[1]_net_1 ), .D(N_1020_1), .Y(sersta64));
    CFG3 #( .INIT(8'hE4) )  \fsmsta_sync_proc.fsmsta_9_am_RNO[2]  (.A(
        un1_fsmsta_nxt_1_sqmuxa_net_1), .B(N_1122), .C(N_1151), .Y(
        N_1128));
    CFG4 #( .INIT(16'h0F08) )  \fsmmod_ns_0[3]  (.A(N_1023), .B(
        \fsmmod[3]_net_1 ), .C(fsmmod5), .D(
        \fsmmod_ns_0_a4_0_4[3]_net_1 ), .Y(\fsmmod_ns[3] ));
    CFG4 #( .INIT(16'hEA00) )  \fsmdet_RNO[6]  (.A(\fsmdet[5]_net_1 ), 
        .B(\fsmdet[6]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_881_i_0));
    CFG4 #( .INIT(16'h78F0) )  
        \framesync_write_proc.framesync_6_enl_bm[3]  (.A(
        \framesync[1]_net_1 ), .B(CO0), .C(\framesync[3]_net_1 ), .D(
        \framesync[2]_net_1 ), .Y(\framesync_6_enl_bm[3] ));
    CFG4 #( .INIT(16'hCCD8) )  \un1_fsmsta_nxt_1[2]  (.A(
        un1_sersta84_1_1_0_net_1), .B(\fsmsta[2]_net_1 ), .C(
        \un1_fsmsta_nxt[2] ), .D(un1_sersta84_1_2_net_1), .Y(
        \un1_fsmsta_nxt_1[2]_net_1 ));
    CFG4 #( .INIT(16'h6626) )  
        \NoName_cnst_2_4_3__NoName_cnst_2_1_0_.m6  (.A(
        \fsmsta[3]_net_1 ), .B(\fsmsta[4]_net_1 ), .C(
        \COREI2C_0_0_SDAO[0] ), .D(SDAInt_net_1), .Y(N_7));
    SLE \serdat[1]  (.D(\serdat_19[1] ), .CLK(GL0_INST), .EN(
        un1_serdat_2_sqmuxa_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\serdat[1]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \un1_SDAInt[0]  (.A(framesync24), .B(
        SDAInt_net_1), .C(\fsmsta[0]_net_1 ), .Y(N_1149));
    CFG4 #( .INIT(16'hCECC) )  un1_sersta60_1 (.A(sersta74_2), .B(
        sersta61), .C(\fsmsta[2]_net_1 ), .D(N_1236_1), .Y(
        un1_sersta60_1_net_1));
    CFG4 #( .INIT(16'h0E00) )  \fsmdet_RNO[3]  (.A(\fsmdet[1]_net_1 ), 
        .B(\fsmdet[6]_net_1 ), .C(SDAInt_net_1), .D(SCLInt_net_1), .Y(
        N_875_i_0));
    CFG4 #( .INIT(16'h2EAA) )  \un1_fsmsta_nxt_2_bm[3]  (.A(
        \NoName_cnst_2[3] ), .B(un1_sersta69_net_1), .C(
        \COREI2C_0_0_SDAO[0] ), .D(framesync24), .Y(
        \un1_fsmsta_nxt_2_bm[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \fsmsync_RNO[1]  (.A(\fsmsync[0]_net_1 ), 
        .B(SCLInt_net_1), .C(N_985), .Y(N_955_i_0));
    CFG4 #( .INIT(16'hF3F2) )  \serdat_write_proc.bsd7_10_iv_1  (.A(
        bsd7_tmp_i_m_1_0), .B(serdat4), .C(\fsmdet[3]_net_1 ), .D(
        \serdat_i_m_0[7] ), .Y(bsd7_10_iv_1));
    CFG3 #( .INIT(8'h48) )  \indelay_4[0]  (.A(\indelay[0]_net_1 ), .B(
        \fsmsync[3]_net_1 ), .C(N_974), .Y(\indelay_4[0]_net_1 ));
    CFG3 #( .INIT(8'hFB) )  \fsmsync_ns_0_o3[0]  (.A(\fsmmod[4]_net_1 )
        , .B(PCLKint_p1_net_1), .C(N_999), .Y(N_972));
    CFG4 #( .INIT(16'hCCCE) )  \fsmmod_ns_0[5]  (.A(N_1048_2), .B(
        N_1047), .C(SDAInt_net_1), .D(N_1031), .Y(\fsmmod_ns[5] ));
    CFG4 #( .INIT(16'h0E00) )  \serdat_write_proc.bsd7_10_iv_1_RNO_0  
        (.A(un1_sersta60_1_net_1), .B(un1_sersta58_1), .C(
        \serdat[7]_net_1 ), .D(bsd7_tmp_7_sn_m6_1_0), .Y(
        \serdat_i_m_0[7] ));
    CFG2 #( .INIT(4'h2) )  PCLKint_p1 (.A(PCLKint_net_1), .B(
        PCLKint_ff_net_1), .Y(PCLKint_p1_net_1));
    SLE \fsmsync[5]  (.D(N_963_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \fsmsync[5]_net_1 ));
    CFG4 #( .INIT(16'hACCC) )  \serdat_write_proc.serdat_19[4]  (.A(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .B(\serdat[3]_net_1 ), .C(
        un1_PSEL), .D(un4_PRDATA), .Y(\serdat_19[4] ));
    CFG4 #( .INIT(16'hF8FA) )  \fsmsync_ns_0_1[0]  (.A(SCLInt_net_1), 
        .B(\fsmsync[4]_net_1 ), .C(N_985), .D(N_980), .Y(
        \fsmsync_ns_0_1[0]_net_1 ));
    CFG4 #( .INIT(16'hFF15) )  
        \framesync_write_proc.framesync_6_enl_am[3]  (.A(framesync10), 
        .B(framesync14), .C(un1_framesync_2), .D(framesync_6_sm0), .Y(
        \framesync_6_enl_am[3] ));
    CFG4 #( .INIT(16'hFFAC) )  ack_RNO (.A(SDAInt_net_1), .B(ack_net_1)
        , .C(un1_serdat_2_sqmuxa_1_net_1), .D(serdat_0_sqmuxa_net_1), 
        .Y(ack_10));
    CFG2 #( .INIT(4'hD) )  \SMBint_filter_proc.SCLI_ff_reg_3[2]  (.A(
        \sercon[6]_net_1 ), .B(\SCLI_ff_reg[1]_net_1 ), .Y(
        \SCLI_ff_reg_3[2] ));
    CFG4 #( .INIT(16'h0010) )  \sercon_write_proc.un1_PRDATA  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(un9_PRDATA_2_0), .D(
        CoreAPB3_0_APBmslave0_PADDR[0]), .Y(un1_PRDATA));
    CFG2 #( .INIT(4'h4) )  nedetect_RNIDG1F (.A(COREI2C_0_0_INT[0]), 
        .B(nedetect_net_1), .Y(bsd7_tmp_7_sn_m6_1_0));
    CFG4 #( .INIT(16'hFFFE) )  \fsmsync_sync_proc.un1_sersta69_1  (.A(
        N_1236), .B(N_1237), .C(sersta77_2), .D(N_1235), .Y(
        un1_sersta69_0));
    CFG4 #( .INIT(16'h0D2F) )  \fsmsta_nxt_3_RNO_0[0]  (.A(
        un1_fsmsta_nxt_2_sn_N_3), .B(un1_framesync24_1_net_1), .C(
        \COREI2C_0_0_SDAO[0] ), .D(N_6), .Y(\un1_fsmsta_nxt_2[0] ));
    CFG4 #( .INIT(16'h1310) )  un1_sersta84_2_1_a6 (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[2]_net_1 ), .C(framesync24), .D(
        N_1020_1), .Y(N_1223));
    CFG2 #( .INIT(4'h1) )  \SDAO_int_write_proc.sersta58_2  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[3]_net_1 ), .Y(sersta74_2));
    SLE \sersta[2]  (.D(\sersta_3[2] ), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sersta[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \fsmsta_comb_proc.fsmsta_nxt19  (.A(
        SDAInt_net_1), .B(\COREI2C_0_0_SDAO[0] ), .Y(fsmsta_nxt19));
    CFG4 #( .INIT(16'hE0EE) )  fsmsta_3_sqmuxa_0_RNIH0MK (.A(
        pedetect_net_1), .B(un1_fsmdet_0), .C(fsmsta13), .D(
        fsmsta_3_sqmuxa_0_net_1), .Y(un1_ens1_pre_1_sqmuxa_i_0));
    CFG4 #( .INIT(16'h0401) )  \sercon_write_proc.un1_framesync_4  (.A(
        \framesync[2]_net_1 ), .B(\framesync[3]_net_1 ), .C(
        \framesync[1]_net_1 ), .D(\framesync[0]_net_1 ), .Y(
        un1_framesync_4));
    CFG4 #( .INIT(16'h0800) )  \fsmsta_sync_proc.fsmsta_9_2_342_i_a3  
        (.A(adrcompen_net_1), .B(un1_framesync24_1_0), .C(sersta64), 
        .D(fsmsta_9_2_342_i_a3_0), .Y(fsmsta_9_2_342_i_a3));
    CFG2 #( .INIT(4'h8) )  \fsmmod_sync_proc.un1_sersta64_0  (.A(
        framesync24), .B(pedetect_net_1), .Y(un1_sersta64_0));
    CFG2 #( .INIT(4'h4) )  nedetect_0_sqmuxa (.A(un1_SCLI_ff_reg), .B(
        SCLInt_net_1), .Y(nedetect_0_sqmuxa_net_1));
    CFG2 #( .INIT(4'h8) )  \SDAO_int_write_proc.sersta75_0  (.A(
        \fsmsta[0]_net_1 ), .B(\fsmsta[4]_net_1 ), .Y(sersta75_0));
    CFG4 #( .INIT(16'hE0A0) )  \indelay_4[2]  (.A(\indelay[2]_net_1 ), 
        .B(\indelay[0]_net_1 ), .C(\fsmsync[3]_net_1 ), .D(
        \indelay[1]_net_1 ), .Y(\indelay_4[2]_net_1 ));
    CFG4 #( .INIT(16'hFFFD) )  \un1_fsmsta_nxt_0_1_iv[2]  (.A(
        \un1_fsmsta_nxt_0_1_iv_1_0[2]_net_1 ), .B(
        \un1_fsmsta_nxt_0_1_iv_1[2]_net_1 ), .C(sersta71), .D(
        un1_sersta60_net_1), .Y(\un1_fsmsta_nxt[2] ));
    CFG2 #( .INIT(4'hE) )  \fsmsta_sync_proc.un1_fsmsta33  (.A(
        un1_fsmmod_1), .B(fsmsta33), .Y(un1_fsmsta33));
    CFG4 #( .INIT(16'h8000) )  \sercon_write_proc.un1_PSEL  (.A(
        un12_PSELi), .B(CoreAPB3_0_APBmslave1_PSELx), .C(
        CoreAPB3_0_APBmslave0_PWRITE), .D(
        CoreAPB3_0_APBmslave0_PENABLE), .Y(un1_PSEL));
    CFG3 #( .INIT(8'hC8) )  \sercon_write_proc.un1_fsmmod_1  (.A(
        \fsmmod[1]_net_1 ), .B(\fsmdet[3]_net_1 ), .C(
        \fsmmod[6]_net_1 ), .Y(un1_fsmmod_1));
    
endmodule


module COREI2C_Z2_layer0(
       COREI2C_0_0_SDAO_i,
       COREI2C_0_0_SCLO_i,
       COREI2C_0_0_INT,
       CoreAPB3_0_APBmslave0_PADDR,
       sersta_m_0,
       sersta_m,
       serdat_m,
       CoreAPB3_0_APBmslave0_PWDATA,
       serdat_4,
       serdat_0,
       sercon_m_6,
       sercon_m_4,
       sercon_m_0,
       \PRDATAi[0]_0 ,
       \PRDATAi[0]_1 ,
       \PRDATAi[0]_2 ,
       \PRDATAi[0]_6 ,
       \PRDATAi[0]_4 ,
       un12_PSELi,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       un9_PRDATA_2_0,
       BIBUF_COREI2C_0_0_SDA_IO_Y,
       BIBUF_COREI2C_0_0_SCL_IO_Y,
       N_528,
       psh_enable_reg1_1_sqmuxa_0,
       un4_PRDATA,
       CoreAPB3_0_APBmslave1_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE
    );
output [0:0] COREI2C_0_0_SDAO_i;
output [0:0] COREI2C_0_0_SCLO_i;
output [0:0] COREI2C_0_0_INT;
input  [8:0] CoreAPB3_0_APBmslave0_PADDR;
output [1:1] sersta_m_0;
output [3:3] sersta_m;
output [6:6] serdat_m;
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output serdat_4;
output serdat_0;
output sercon_m_6;
output sercon_m_4;
output sercon_m_0;
output \PRDATAi[0]_0 ;
output \PRDATAi[0]_1 ;
output \PRDATAi[0]_2 ;
output \PRDATAi[0]_6 ;
output \PRDATAi[0]_4 ;
output un12_PSELi;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output un9_PRDATA_2_0;
input  BIBUF_COREI2C_0_0_SDA_IO_Y;
input  BIBUF_COREI2C_0_0_SCL_IO_Y;
input  N_528;
input  psh_enable_reg1_1_sqmuxa_0;
output un4_PRDATA;
input  CoreAPB3_0_APBmslave1_PSELx;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    COREI2CREAL_Z3_layer0 \I2C_NUM_GENERATION[0].ui2c  (
        .COREI2C_0_0_SDAO_i({COREI2C_0_0_SDAO_i[0]}), 
        .COREI2C_0_0_SCLO_i({COREI2C_0_0_SCLO_i[0]}), .COREI2C_0_0_INT({
        COREI2C_0_0_INT[0]}), .CoreAPB3_0_APBmslave0_PADDR({
        CoreAPB3_0_APBmslave0_PADDR[4], CoreAPB3_0_APBmslave0_PADDR[3], 
        CoreAPB3_0_APBmslave0_PADDR[2], CoreAPB3_0_APBmslave0_PADDR[1], 
        CoreAPB3_0_APBmslave0_PADDR[0]}), .sersta_m_0({sersta_m_0[1]}), 
        .serdat_m({serdat_m[6]}), .CoreAPB3_0_APBmslave0_PWDATA({
        CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .serdat_4(serdat_4), 
        .serdat_0(serdat_0), .sersta_m_3(sersta_m[3]), .sercon_m_6(
        sercon_m_6), .sercon_m_4(sercon_m_4), .sercon_m_0(sercon_m_0), 
        .\PRDATAi[0]_0 (\PRDATAi[0]_0 ), .\PRDATAi[0]_1 (
        \PRDATAi[0]_1 ), .\PRDATAi[0]_2 (\PRDATAi[0]_2 ), 
        .\PRDATAi[0]_6 (\PRDATAi[0]_6 ), .\PRDATAi[0]_4 (
        \PRDATAi[0]_4 ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .un9_PRDATA_2_0(un9_PRDATA_2_0), .BIBUF_COREI2C_0_0_SDA_IO_Y(
        BIBUF_COREI2C_0_0_SDA_IO_Y), .BIBUF_COREI2C_0_0_SCL_IO_Y(
        BIBUF_COREI2C_0_0_SCL_IO_Y), .N_528(N_528), 
        .psh_enable_reg1_1_sqmuxa_0(psh_enable_reg1_1_sqmuxa_0), 
        .un4_PRDATA(un4_PRDATA), .un12_PSELi(un12_PSELi), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0001) )  \I2C_NUM_PSELi_GEN[0].un12_PSELi  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[8]), .D(
        CoreAPB3_0_APBmslave0_PADDR[6]), .Y(un12_PSELi));
    
endmodule


module CoreResetP_Z6_layer0(
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       SYSRESET_POR,
       mss_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N
    );
output MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  SYSRESET_POR;
input  mss_sb_MSS_TMP_0_MSS_RESET_N_M2F;
input  mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N;

    wire MSS_HPMS_READY_int_net_1, mss_ready_select_net_1, VCC_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        GND_net_1, mss_ready_state_net_1, RESET_N_M2F_clk_base_net_1, 
        POWER_ON_RESET_N_q1_net_1, RESET_N_M2F_q1_net_1, 
        FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, MSS_HPMS_READY_int_4_net_1;
    
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(RESET_N_M2F_clk_base_net_1));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_clk_base_net_1));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        mss_ready_select4_net_1), .ALn(POWER_ON_RESET_N_clk_base_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(mss_ready_select_net_1));
    CLKINT MSS_HPMS_READY_int_RNI5CTC_inst_1 (.A(
        MSS_HPMS_READY_int_net_1), .Y(MSS_HPMS_READY_int_RNI5CTC));
    GND GND (.Y(GND_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        RESET_N_M2F_clk_base_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_q1_net_1));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_q1_net_1));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Rx_async_1s_0s_1s_2s(
       rx_byte,
       controlReg2,
       clear_parity_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       Echo_control_0_TX,
       CoreUARTapb_2_0_PARITY_ERR,
       stop_strobe,
       CoreUARTapb_2_0_FRAMING_ERR,
       clear_parity_en,
       fifo_write,
       rx_idle
    );
output [7:0] rx_byte;
input  [2:0] controlReg2;
input  clear_parity_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  baud_clock;
input  Echo_control_0_TX;
output CoreUARTapb_2_0_PARITY_ERR;
output stop_strobe;
output CoreUARTapb_2_0_FRAMING_ERR;
output clear_parity_en;
output fifo_write;
output rx_idle;

    wire clear_parity_reg_i_0, \rx_bit_cnt[0]_net_1 , VCC_net_1, 
        N_326_i_0, GND_net_1, \rx_bit_cnt[1]_net_1 , N_325_i_0, 
        \rx_bit_cnt[2]_net_1 , N_324_i_0, \rx_bit_cnt[3]_net_1 , 
        N_323_i_0, \samples[1]_net_1 , \samples[2]_net_1 , 
        \rx_shift[0]_net_1 , \rx_shift_11[0] , 
        un1_samples7_1_0_0_net_1, \rx_shift[1]_net_1 , 
        \rx_shift_11[1] , \rx_shift[2]_net_1 , \rx_shift_11[2] , 
        \rx_shift[3]_net_1 , \rx_shift_11[3] , \rx_shift[4]_net_1 , 
        \rx_shift_11[4] , \rx_shift[5]_net_1 , \rx_shift_11[5] , 
        \rx_shift[6]_net_1 , N_322_i_0, \rx_shift[7]_net_1 , N_283_i_0, 
        \rx_shift[8]_net_1 , N_282_i_0, \receive_count[0]_net_1 , 
        N_287_i_0, \receive_count[1]_net_1 , N_286_i_0, 
        \receive_count[2]_net_1 , N_285_i_0, \receive_count[3]_net_1 , 
        N_284_i_0, clear_parity_en_9, N_288_i_0, \samples[0]_net_1 , 
        N_310, parity_err_1_sqmuxa_i_0_net_1, rx_parity_calc_net_1, 
        N_321_i_0, framing_error_int_net_1, framing_error_int_0_sqmuxa, 
        framing_error_int_2_sqmuxa, framing_error_1_sqmuxa_i_0_net_1, 
        \rx_state[1]_net_1 , N_233_i_0, \rx_state[0]_net_1 , 
        \rx_state_ns[0] , clear_parity_en_9_i_0, N_331, N_350, N_124, 
        rx_state19_NE_1, rx_state19_li, N_332, 
        framing_error_int_0_sqmuxa_0_a2_0_net_1, 
        \rx_state_ns_i_0_a2_0_0[1] , N_357_1, 
        parity_err_1_sqmuxa_i_a2_0_1_net_1, 
        parity_err_1_sqmuxa_i_a2_2_net_1, N_293, \rx_shift_11_i_0[7] , 
        N_126, N_329, N_174, N_314, N_77, 
        parity_err_1_sqmuxa_i_0_0_net_1, N_58;
    
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[2]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  \rcv_cnt.receive_count_3_i_a2[0]  (.A(
        \receive_count[1]_net_1 ), .B(rx_idle), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[3]_net_1 ), .Y(
        N_126));
    CFG3 #( .INIT(8'h06) )  \receive_shift.rx_shift_11_i_a2[7]  (.A(
        controlReg2[0]), .B(controlReg2[1]), .C(N_329), .Y(N_314));
    CFG2 #( .INIT(4'h8) )  framing_error_int_0_sqmuxa_0_a2_1 (.A(
        \rx_state[1]_net_1 ), .B(\receive_count[2]_net_1 ), .Y(
        \rx_state_ns_i_0_a2_0_0[1] ));
    CFG2 #( .INIT(4'h4) )  framing_error_int_0_sqmuxa_0_a2_0 (.A(
        \receive_count[0]_net_1 ), .B(\receive_count[1]_net_1 ), .Y(
        framing_error_int_0_sqmuxa_0_a2_0_net_1));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[0]));
    CFG4 #( .INIT(16'h0004) )  \rcv_cnt.receive_count_3_i_a2_0[3]  (.A(
        \receive_count[0]_net_1 ), .B(rx_idle), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_174));
    SLE \receive_count[1]  (.D(N_286_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[1]_net_1 ));
    SLE \rx_shift[7]  (.D(N_283_i_0), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[7]_net_1 ));
    CFG3 #( .INIT(8'hBA) )  \receive_shift.rx_shift_11_i_0[7]  (.A(
        rx_idle), .B(\rx_shift[8]_net_1 ), .C(N_357_1), .Y(
        \rx_shift_11_i_0[7] ));
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[0]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \receive_shift.rx_shift_11_i_o2[6]  (.A(
        controlReg2[1]), .B(controlReg2[0]), .Y(N_332));
    CFG1 #( .INIT(2'h1) )  framing_error_RNO (.A(clear_parity_reg), .Y(
        clear_parity_reg_i_0));
    CFG3 #( .INIT(8'h02) )  parity_err_1_sqmuxa_i_a2_0_1 (.A(
        controlReg2[1]), .B(\rx_bit_cnt[3]_net_1 ), .C(controlReg2[0]), 
        .Y(parity_err_1_sqmuxa_i_a2_0_1_net_1));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[0]  (.A(rx_idle), 
        .B(\rx_shift[1]_net_1 ), .Y(\rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(N_284_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[3]_net_1 ));
    CFG4 #( .INIT(16'h0096) )  
        \make_parity_err.parity_err_12_iv_0_111_a2_0_a2  (.A(
        controlReg2[2]), .B(rx_parity_calc_net_1), .C(N_329), .D(
        clear_parity_reg), .Y(N_310));
    VCC VCC (.Y(VCC_net_1));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[4]));
    CFG3 #( .INIT(8'h7F) )  \rcv_cnt.receive_count_3_i_o2_0[2]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(N_293));
    CFG4 #( .INIT(16'h333B) )  un1_samples7_1_0_0 (.A(baud_clock), .B(
        N_331), .C(\rx_state[1]_net_1 ), .D(\rx_state[0]_net_1 ), .Y(
        un1_samples7_1_0_0_net_1));
    SLE rx_parity_calc (.D(N_321_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_parity_calc_net_1));
    SLE \rx_bit_cnt[2]  (.D(N_324_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[2]_net_1 ));
    SLE \rx_bit_cnt[1]  (.D(N_325_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[1]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \rx_state_RNI1CK2[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(rx_idle));
    CFG3 #( .INIT(8'h21) )  rx_parity_calc_RNO (.A(
        rx_parity_calc_net_1), .B(\rx_state[1]_net_1 ), .C(N_77), .Y(
        N_321_i_0));
    CFG3 #( .INIT(8'h09) )  \rx_bit_cnt_RNO[0]  (.A(N_331), .B(
        \rx_bit_cnt[0]_net_1 ), .C(N_350), .Y(N_326_i_0));
    CFG4 #( .INIT(16'h1230) )  \receive_count_RNO[2]  (.A(
        \receive_count[0]_net_1 ), .B(N_124), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_285_i_0));
    CFG4 #( .INIT(16'h0240) )  \rcv_sm.rx_state19_NE_1  (.A(
        \rx_bit_cnt[1]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(N_332), 
        .D(\rx_bit_cnt[2]_net_1 ), .Y(rx_state19_NE_1));
    SLE stop_strobe_inst_1 (.D(framing_error_int_2_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG4 #( .INIT(16'h3022) )  \rx_shift_RNO[6]  (.A(N_329), .B(
        rx_idle), .C(\rx_shift[7]_net_1 ), .D(N_332), .Y(N_322_i_0));
    CFG4 #( .INIT(16'h00CE) )  \rx_state_RNO[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .C(
        rx_state19_li), .D(framing_error_int_2_sqmuxa), .Y(N_233_i_0));
    CFG3 #( .INIT(8'h09) )  \rx_bit_cnt_RNO[2]  (.A(N_58), .B(
        \rx_bit_cnt[2]_net_1 ), .C(N_350), .Y(N_324_i_0));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[1]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[2]  (.A(rx_idle), 
        .B(\rx_shift[3]_net_1 ), .Y(\rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(N_285_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[2]_net_1 ));
    SLE clear_parity_en_1 (.D(clear_parity_en_9), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_en));
    CFG4 #( .INIT(16'hF2F0) )  parity_err_1_sqmuxa_i_0_0 (.A(
        parity_err_1_sqmuxa_i_a2_2_net_1), .B(N_331), .C(
        clear_parity_reg), .D(N_357_1), .Y(
        parity_err_1_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'hBAAA) )  parity_err_1_sqmuxa_i_0 (.A(
        parity_err_1_sqmuxa_i_0_0_net_1), .B(N_58), .C(
        \rx_bit_cnt[2]_net_1 ), .D(parity_err_1_sqmuxa_i_a2_0_1_net_1), 
        .Y(parity_err_1_sqmuxa_i_0_net_1));
    SLE \rx_state[1]  (.D(N_233_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    CFG4 #( .INIT(16'h000E) )  \rx_shift_RNO[7]  (.A(
        \rx_shift[7]_net_1 ), .B(N_332), .C(\rx_shift_11_i_0[7] ), .D(
        N_314), .Y(N_283_i_0));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[6]));
    CFG3 #( .INIT(8'h12) )  \receive_count_RNO[1]  (.A(
        \receive_count[0]_net_1 ), .B(N_124), .C(
        \receive_count[1]_net_1 ), .Y(N_286_i_0));
    GND GND (.Y(GND_net_1));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[3]  (.A(rx_idle), 
        .B(\rx_shift[4]_net_1 ), .Y(\rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(N_288_i_0), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[7]));
    CFG4 #( .INIT(16'h7BB7) )  \rcv_sm.rx_state19_NE  (.A(
        controlReg2[1]), .B(rx_state19_NE_1), .C(\rx_bit_cnt[0]_net_1 )
        , .D(controlReg2[0]), .Y(rx_state19_li));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[3]));
    CFG3 #( .INIT(8'h40) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_0_a2  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9));
    CFG4 #( .INIT(16'h1001) )  \receive_count_RNO[3]  (.A(N_174), .B(
        N_124), .C(\receive_count[3]_net_1 ), .D(N_293), .Y(N_284_i_0));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[2]));
    CFG3 #( .INIT(8'hE8) )  \rx_filtered.m3_0_o2  (.A(
        \samples[1]_net_1 ), .B(\samples[0]_net_1 ), .C(
        \samples[2]_net_1 ), .Y(N_329));
    CFG3 #( .INIT(8'h01) )  \receive_count_RNO[0]  (.A(N_124), .B(
        \receive_count[0]_net_1 ), .C(N_126), .Y(N_287_i_0));
    SLE parity_err (.D(N_310), .CLK(GL0_INST), .EN(
        parity_err_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(CoreUARTapb_2_0_PARITY_ERR)
        );
    SLE \rx_shift[6]  (.D(N_322_i_0), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[6]_net_1 ));
    CFG3 #( .INIT(8'h04) )  \receive_shift.rx_bit_cnt_4_i_a2[3]  (.A(
        \rx_state[0]_net_1 ), .B(baud_clock), .C(\rx_state[1]_net_1 ), 
        .Y(N_350));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[4]  (.A(rx_idle), 
        .B(\rx_shift[5]_net_1 ), .Y(\rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[3]_net_1 ));
    SLE framing_error_int (.D(framing_error_int_0_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(framing_error_int_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \rx_state_ns_0_0[0]  (.A(N_174), .B(
        rx_state19_li), .C(\rx_state[0]_net_1 ), .D(
        \receive_count[3]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \samples[2]  (.D(Echo_control_0_TX), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    SLE \receive_count[0]  (.D(N_287_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[5]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[5]  (.A(rx_idle), 
        .B(\rx_shift[6]_net_1 ), .Y(\rx_shift_11[5] ));
    CFG4 #( .INIT(16'h8000) )  \rx_state_ns_i_0_a2_0[1]  (.A(
        \receive_count[0]_net_1 ), .B(\rx_state_ns_i_0_a2_0_0[1] ), .C(
        \receive_count[3]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        framing_error_int_2_sqmuxa));
    CFG4 #( .INIT(16'h0800) )  framing_error_int_0_sqmuxa_0_a2 (.A(
        framing_error_int_0_sqmuxa_0_a2_0_net_1), .B(
        \receive_count[3]_net_1 ), .C(N_329), .D(
        \rx_state_ns_i_0_a2_0_0[1] ), .Y(framing_error_int_0_sqmuxa));
    CFG3 #( .INIT(8'hDF) )  \receive_shift.rx_bit_cnt_4_i_o2[2]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(N_331), .C(\rx_bit_cnt[1]_net_1 ), 
        .Y(N_58));
    CFG4 #( .INIT(16'h0002) )  parity_err_1_sqmuxa_i_a2_2 (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        \rx_bit_cnt[2]_net_1 ), .D(\rx_bit_cnt[0]_net_1 ), .Y(
        parity_err_1_sqmuxa_i_a2_2_net_1));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[5]_net_1 ));
    CFG4 #( .INIT(16'hE800) )  \rcv_cnt.receive_count_3_i_a2[3]  (.A(
        \samples[0]_net_1 ), .B(\samples[1]_net_1 ), .C(
        \samples[2]_net_1 ), .D(rx_idle), .Y(N_124));
    SLE \rx_bit_cnt[0]  (.D(N_326_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[0]_net_1 ));
    SLE \rx_shift[8]  (.D(N_282_i_0), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rx_shift[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[1]  (.A(rx_idle), 
        .B(\rx_shift[2]_net_1 ), .Y(\rx_shift_11[1] ));
    CFG3 #( .INIT(8'hDF) )  \receive_shift.rx_bit_cnt_4_i_o2[0]  (.A(
        baud_clock), .B(N_293), .C(\receive_count[3]_net_1 ), .Y(N_331)
        );
    CFG3 #( .INIT(8'hBF) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_0_a2_i  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9_i_0));
    SLE framing_error (.D(clear_parity_reg_i_0), .CLK(GL0_INST), .EN(
        framing_error_1_sqmuxa_i_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_0_FRAMING_ERR));
    CFG4 #( .INIT(16'hFF7F) )  \rx_par_calc.rx_parity_calc_4_u_i_o2  (
        .A(controlReg2[1]), .B(\receive_count[3]_net_1 ), .C(N_329), 
        .D(N_293), .Y(N_77));
    CFG3 #( .INIT(8'hEC) )  framing_error_1_sqmuxa_i_0 (.A(
        framing_error_int_net_1), .B(clear_parity_reg), .C(baud_clock), 
        .Y(framing_error_1_sqmuxa_i_0_net_1));
    CFG4 #( .INIT(16'h2230) )  \rx_shift_RNO[8]  (.A(N_329), .B(
        rx_idle), .C(\rx_shift[8]_net_1 ), .D(N_357_1), .Y(N_282_i_0));
    CFG2 #( .INIT(4'h8) )  \rx_byte_RNO[7]  (.A(controlReg2[0]), .B(
        \rx_shift[7]_net_1 ), .Y(N_288_i_0));
    CFG4 #( .INIT(16'h0A06) )  \rx_bit_cnt_RNO[3]  (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(N_350), 
        .D(N_58), .Y(N_323_i_0));
    CFG2 #( .INIT(4'h8) )  parity_err_1_sqmuxa_i_a2_1 (.A(
        controlReg2[1]), .B(controlReg2[0]), .Y(N_357_1));
    SLE \rx_bit_cnt[3]  (.D(N_323_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h0A06) )  \rx_bit_cnt_RNO[1]  (.A(
        \rx_bit_cnt[1]_net_1 ), .B(\rx_bit_cnt[0]_net_1 ), .C(N_350), 
        .D(N_331), .Y(N_325_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_0_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] tx_hold_reg;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), .C_WEN(
        INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), 
        .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_ctrl_128(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_3704_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, \counter[0]_net_1 , 
        VCC_net_1, un1_counter_cry_0_Y_2, GND_net_1, 
        \counter[1]_net_1 , un1_counter_cry_1_0_S_1, 
        \counter[2]_net_1 , un1_counter_cry_2_0_S_1, 
        \counter[3]_net_1 , un1_counter_cry_3_0_S_1, 
        \counter[4]_net_1 , un1_counter_cry_4_0_S_1, 
        \counter[5]_net_1 , un1_counter_cry_5_0_S_1, 
        \counter[6]_net_1 , un1_counter_s_6_S_1, \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \data_out_0[0] , 
        \data_out_0[1] , \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_312_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_313_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        empty_4_net_1, full_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_313_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_2_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[2]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S_1), .Y(), .FCO(
        un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[3]));
    CFG4 #( .INIT(16'h7FFF) )  full_4_RNIGLBA (.A(\counter[0]_net_1 ), 
        .B(full_4_net_1), .C(\counter[6]_net_1 ), .D(
        \counter[4]_net_1 ), .Y(fifo_full_tx_i_0));
    SLE \counter[6]  (.D(un1_counter_s_6_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_4_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[4]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S_1), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_312_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIHRB7 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[6]));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_3_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[3]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S_1), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_tx), .C(fifo_write_tx), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_2), 
        .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[4]_net_1 ), 
        .Y(fifo_empty_tx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_3704_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_312 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_312_FCO));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_313 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_313_FCO));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_1_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_1), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    CFG1 #( .INIT(2'h1) )  N_3704_i_0 (.A(fifo_write_tx), .Y(
        N_3704_i_0_net_1));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_5_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[5]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S_1), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_0_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg({
        tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], 
        tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]})
        , .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_tx(fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(\counter[6]_net_1 ), 
        .FCI(un1_counter_cry_5), .S(un1_counter_s_6_S_1), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_256x8(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_0_fifo_ctrl_128 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.tx_dout_reg({
        tx_dout_reg[7], tx_dout_reg[6], tx_dout_reg[5], tx_dout_reg[4], 
        tx_dout_reg[3], tx_dout_reg[2], tx_dout_reg[1], tx_dout_reg[0]})
        , .tx_hold_reg({tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], 
        tx_hold_reg[4], tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], 
        tx_hold_reg[0]}), .fifo_write_tx(fifo_write_tx), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       controlReg2,
       fifo_read_tx,
       fifo_read_tx_i_0,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_289,
       mss_sb_0_TX,
       CoreUARTapb_2_0_TXRDY,
       fifo_full_tx_i_0,
       xmit_clock,
       baud_clock,
       fifo_empty_tx
    );
input  [7:0] tx_dout_reg;
input  [2:0] controlReg2;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_289;
output mss_sb_0_TX;
output CoreUARTapb_2_0_TXRDY;
input  fifo_full_tx_i_0;
input  xmit_clock;
input  baud_clock;
input  fifo_empty_tx;

    wire \tx_byte[4]_net_1 , VCC_net_1, N_133_i_0, GND_net_1, 
        \tx_byte[5]_net_1 , \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_122_i_0, \xmit_bit_sel[2]_net_1 , 
        N_124_i_0, \xmit_bit_sel[3]_net_1 , N_126_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , \tx_byte[2]_net_1 , 
        \tx_byte[3]_net_1 , tx_parity_net_1, tx_parity_5, 
        un1_tx_parity_1_sqmuxa_0_0_net_1, tx_4_iv_i_0, N_144_i_0, 
        \xmit_state_ns_i_0[6] , \xmit_state[6]_net_1 , 
        \xmit_state_ns[6] , \xmit_state[0]_net_1 , \xmit_state_ns[0] , 
        \xmit_state[1]_net_1 , \xmit_state[2]_net_1 , 
        \xmit_state_ns[2]_net_1 , \xmit_state[3]_net_1 , N_112_i_0, 
        \xmit_state[4]_net_1 , \xmit_state_ns[4] , 
        \xmit_state[5]_net_1 , \xmit_state_ns[5] , N_176, 
        tx_2_u_i_m2_am_1_1, tx_2_u_i_m2_am, tx_2_u_i_m2_bm_1_1, 
        tx_2_u_i_m2_bm, N_473, N_82, N_80_i, N_130, N_173, N_132;
    
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(
        tx_2_u_i_m2_bm_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_bm));
    SLE tx_parity (.D(tx_parity_5), .CLK(GL0_INST), .EN(
        un1_tx_parity_1_sqmuxa_0_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_parity_net_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_0_TXRDY));
    CFG4 #( .INIT(16'h8000) )  un1_tx_parity_1_sqmuxa_0_0_a2 (.A(
        \xmit_state[3]_net_1 ), .B(xmit_clock), .C(baud_clock), .D(
        controlReg2[1]), .Y(N_176));
    CFG3 #( .INIT(8'hD8) )  \xmit_sel.tx_2_u_i_m2_ns  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(tx_2_u_i_m2_bm), .C(
        tx_2_u_i_m2_am), .Y(N_473));
    SLE \xmit_state[3]  (.D(N_112_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[3]_net_1 ));
    CFG4 #( .INIT(16'h0501) )  \xmit_sel.tx_4_iv_i  (.A(
        \xmit_state[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_130), 
        .D(N_473), .Y(tx_4_iv_i_0));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[0]_net_1 ));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNI169 (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    CFG4 #( .INIT(16'hFCFA) )  \xmit_state_ns_0[5]  (.A(
        \xmit_state[5]_net_1 ), .B(\xmit_state[4]_net_1 ), .C(N_132), 
        .D(N_289), .Y(\xmit_state_ns[5] ));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3_0_a2[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[0]_net_1 ), .B(\xmit_bit_sel[1]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_122_i_0));
    CFG2 #( .INIT(4'h7) )  \xmit_cnt.xmit_bit_sel_3_i_0_o2[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(N_82)
        );
    CFG2 #( .INIT(4'h8) )  \xmit_state_RNI7UIQ[2]  (.A(N_289), .B(
        \xmit_state[2]_net_1 ), .Y(N_133_i_0));
    VCC VCC (.Y(VCC_net_1));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[5]_net_1 ));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_bm_1_1));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[5]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_state_RNI0IIN1[1]  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(N_289), 
        .D(\xmit_state[6]_net_1 ), .Y(N_144_i_0));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(N_289), 
        .Y(\xmit_state_ns[2]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \xmit_state_ns_0_a2[5]  (.A(
        controlReg2[1]), .B(\xmit_state[3]_net_1 ), .C(N_289), .D(
        N_173), .Y(N_132));
    CFG4 #( .INIT(16'h0200) )  \xmit_state_ns_0_a2_0[5]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(N_80_i), .C(
        \xmit_bit_sel[3]_net_1 ), .D(\xmit_bit_sel[2]_net_1 ), .Y(
        N_173));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_126_i_0), .CLK(GL0_INST), .EN(N_289), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[3]_net_1 ));
    CFG3 #( .INIT(8'h82) )  \xmit_sel.tx_4_iv_0_a2_0  (.A(
        \xmit_state[4]_net_1 ), .B(controlReg2[2]), .C(tx_parity_net_1)
        , .Y(N_130));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns_0[0]  (.A(fifo_empty_tx), 
        .B(N_289), .C(\xmit_state[5]_net_1 ), .D(\xmit_state[0]_net_1 )
        , .Y(\xmit_state_ns[0] ));
    SLE \xmit_bit_sel[2]  (.D(N_124_i_0), .CLK(GL0_INST), .EN(N_289), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'hB) )  fifo_read_en0_1_i_a3_0_a2_i (.A(
        fifo_empty_tx), .B(\xmit_state[0]_net_1 ), .Y(
        \xmit_state_ns_i_0[6] ));
    SLE tx (.D(tx_4_iv_i_0), .CLK(GL0_INST), .EN(N_144_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(mss_sb_0_TX));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[3]_net_1 ));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[7]_net_1 ));
    CFG4 #( .INIT(16'hAECC) )  \xmit_state_RNO[3]  (.A(
        \xmit_state[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_173), 
        .D(N_289), .Y(N_112_i_0));
    CFG3 #( .INIT(8'h12) )  \xmit_par_calc.tx_parity_5  (.A(
        tx_parity_net_1), .B(\xmit_state[5]_net_1 ), .C(N_473), .Y(
        tx_parity_5));
    CFG3 #( .INIT(8'h84) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_82), 
        .Y(N_124_i_0));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_tx_parity_1_sqmuxa_0_0 (.A(N_176), .B(
        \xmit_state[5]_net_1 ), .Y(un1_tx_parity_1_sqmuxa_0_0_net_1));
    SLE \xmit_bit_sel[1]  (.D(N_122_i_0), .CLK(GL0_INST), .EN(N_289), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  fifo_read_en0_1_i_a3_0_a2 (.A(fifo_empty_tx)
        , .B(\xmit_state[0]_net_1 ), .Y(\xmit_state_ns[6] ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[1]_net_1 ));
    CFG4 #( .INIT(16'hC0EA) )  \xmit_state_ns_0[4]  (.A(
        \xmit_state[4]_net_1 ), .B(N_176), .C(N_173), .D(N_289), .Y(
        \xmit_state_ns[4] ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(GL0_INST), 
        .EN(N_289), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[2]_net_1 ));
    SLE fifo_read_en0 (.D(\xmit_state_ns_i_0[6] ), .CLK(GL0_INST), .EN(
        N_144_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    CFG2 #( .INIT(4'h6) )  \xmit_state_ns_0_x2[5]  (.A(controlReg2[0]), 
        .B(\xmit_bit_sel[0]_net_1 ), .Y(N_80_i));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[1]_net_1 ));
    SLE \xmit_state[4]  (.D(\xmit_state_ns[4] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[4]_net_1 ));
    CFG4 #( .INIT(16'hC600) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_bit_sel[3]_net_1 ), .C(N_82)
        , .D(\xmit_state[3]_net_1 ), .Y(N_126_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_am_1_1));
    SLE \xmit_state[6]  (.D(\xmit_state_ns[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[6]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(
        tx_2_u_i_m2_am_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_am));
    
endmodule


module mss_sb_CoreUARTapb_2_0_Clock_gen_0s(
       controlReg1,
       controlReg2,
       xmit_clock,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       N_289
    );
input  [7:0] controlReg1;
input  [7:3] controlReg2;
output xmit_clock;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output baud_clock;
output N_289;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNIQ6LQ_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI89KCK[11]  (.A(
        VCC_net_1), .B(controlReg2[6]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[11] ), .FCI(\baud_cntr_cry[10] ), .S(
        \baud_cntr_s[11] ), .Y(), .FCO(\baud_cntr_cry[11] ));
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIRMIG2[0]  (.A(
        VCC_net_1), .B(controlReg1[0]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[0] ), .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), 
        .Y(), .FCO(\baud_cntr_cry[0] ));
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[1] ));
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[3] ));
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[3]_net_1 ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[9] ));
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNIQ6LQ_Y), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(baud_clock));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIQ03AE[7]  (.A(
        VCC_net_1), .B(controlReg1[7]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[7] ), .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] )
        , .Y(), .FCO(\baud_cntr_cry[7] ));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[7] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[5] ));
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIAJBI7[3]  (.A(
        VCC_net_1), .B(controlReg1[3]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[3] ), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] )
        , .Y(), .FCO(\baud_cntr_cry[3] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI3TDS5[2]  (.A(
        VCC_net_1), .B(controlReg1[2]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[2] ), .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] )
        , .Y(), .FCO(\baud_cntr_cry[2] ));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[0] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIB25KC[6]  (.A(
        VCC_net_1), .B(controlReg1[6]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[6] ), .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] )
        , .Y(), .FCO(\baud_cntr_cry[6] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIJB989[4]  (.A(
        VCC_net_1), .B(controlReg1[4]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[4] ), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] )
        , .Y(), .FCO(\baud_cntr_cry[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIU8G64[1]  (.A(
        VCC_net_1), .B(controlReg1[1]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[1] ), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] )
        , .Y(), .FCO(\baud_cntr_cry[1] ));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIMV4OH[9]  (.A(
        VCC_net_1), .B(controlReg2[4]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[9] ), .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] )
        , .Y(), .FCO(\baud_cntr_cry[9] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[6] ));
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        xmit_clock));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNIQ6LQ  (.A(baud_cntr8_8)
        , .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(baud_cntr8_7), .FCI(
        VCC_net_1), .S(), .Y(baud_cntr8_1_RNIQ6LQ_Y), .FCO(
        baud_cntr_cry_cy));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIU57UA[5]  (.A(
        VCC_net_1), .B(controlReg1[5]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[5] ), .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] )
        , .Y(), .FCO(\baud_cntr_cry[5] ));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h44700) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(controlReg2[7]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[12] ), .FCI(\baud_cntr_cry[11] ), .S(
        \baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[1]_net_1 ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI7V31G[8]  (.A(
        VCC_net_1), .B(controlReg2[3]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[8] ), .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] )
        , .Y(), .FCO(\baud_cntr_cry[8] ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[2] ));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIEJC2J[10]  (.A(
        VCC_net_1), .B(controlReg2[5]), .C(baud_cntr8_1_RNIQ6LQ_Y), .D(
        \baud_cntr[10] ), .FCI(\baud_cntr_cry[9] ), .S(
        \baud_cntr_s[10] ), .Y(), .FCO(\baud_cntr_cry[10] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    CFG2 #( .INIT(4'h8) )  xmit_pulse_i_1_o2 (.A(baud_clock), .B(
        xmit_clock), .Y(N_289));
    
endmodule


module mss_sb_CoreUARTapb_2_0_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte_in,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       N_347_i_0
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte_in;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  N_347_i_0;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte_in[7], rx_byte_in[6], 
        rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], 
        rx_byte_in[1], rx_byte_in[0]}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(N_347_i_0), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_ctrl_128_0(
       rx_dout,
       rx_state,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_write_rx_1_i_a2_0_a2,
       N_347_i_0,
       rx_dout_reg_empty,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [1:0] rx_state;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_write_rx_1_i_a2_0_a2;
input  N_347_i_0;
input  rx_dout_reg_empty;
output fifo_empty_rx;
output fifo_full_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[1]_net_1 , VCC_net_1, 
        un1_counter_cry_1_0_S_2, GND_net_1, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_2, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S_2, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_2, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_2, \counter[6]_net_1 , 
        un1_counter_s_6_S_2, \counter[0]_net_1 , un1_counter_cry_0_Y_1, 
        \data_out_0[0] , \data_out_0[1] , \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , empty_RNI0RU31_net_1, 
        \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , N_295_i_0, 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_314_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_315_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_4_net_1, empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_315_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIG41E (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_2_0 (.A(N_295_i_0), .B(
        N_347_i_0), .C(\counter[2]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S_2), .Y(), .FCO(
        un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(empty_RNI0RU31_net_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_4_0 (.A(N_295_i_0), .B(
        N_347_i_0), .C(\counter[4]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S_2), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_314_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_write_rx_1_i_a2_0_a2), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_2), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_3_0 (.A(N_295_i_0), .B(
        N_347_i_0), .C(\counter[3]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S_2), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_314 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_314_FCO));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(empty_RNI0RU31_net_1), .C(N_347_i_0), 
        .D(GND_net_1), .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_1)
        , .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_empty_rx));
    CFG4 #( .INIT(16'h0004) )  empty_RNI0RU31_0 (.A(rx_state[1]), .B(
        rx_dout_reg_empty), .C(fifo_empty_rx), .D(rx_state[0]), .Y(
        N_295_i_0));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_write_rx_1_i_a2_0_a2), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_315 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_315_FCO));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_1_0 (.A(N_295_i_0), .B(
        N_347_i_0), .C(\counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_2), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[1]));
    CFG4 #( .INIT(16'h8000) )  full (.A(\counter[0]_net_1 ), .B(
        full_4_net_1), .C(\counter[3]_net_1 ), .D(\counter[1]_net_1 ), 
        .Y(fifo_full_rx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_5_0 (.A(N_295_i_0), .B(
        N_347_i_0), .C(\counter[5]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S_2), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_295_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_0_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte_in({
        rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], 
        rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .N_347_i_0(N_347_i_0));
    CFG4 #( .INIT(16'hFFFB) )  empty_RNI0RU31 (.A(rx_state[1]), .B(
        rx_dout_reg_empty), .C(fifo_empty_rx), .D(rx_state[0]), .Y(
        empty_RNI0RU31_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h46A00) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        \counter[6]_net_1 ), .C(N_295_i_0), .D(N_347_i_0), .FCI(
        un1_counter_cry_5), .S(un1_counter_s_6_S_2), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_1), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[2]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_0_fifo_256x8_0(
       rx_dout,
       rx_state,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_write_rx_1_i_a2_0_a2,
       N_347_i_0,
       rx_dout_reg_empty,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [1:0] rx_state;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_write_rx_1_i_a2_0_a2;
input  N_347_i_0;
input  rx_dout_reg_empty;
output fifo_empty_rx;
output fifo_full_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_0_fifo_ctrl_128_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_state({rx_state[1], rx_state[0]})
        , .rx_byte_in({rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], 
        rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], 
        rx_byte_in[0]}), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .fifo_write_rx_1_i_a2_0_a2(fifo_write_rx_1_i_a2_0_a2), 
        .N_347_i_0(N_347_i_0), .rx_dout_reg_empty(rx_dout_reg_empty), 
        .fifo_empty_rx(fifo_empty_rx), .fifo_full_rx(fifo_full_rx));
    
endmodule


module mss_sb_CoreUARTapb_2_0_COREUART_1s_1s_0s_15s_0s(
       CoreAPB3_0_APBmslave0_PWDATA,
       data_out,
       CoreAPB3_0_APBmslave0_PADDR,
       controlReg1,
       controlReg2,
       rx_dout_reg_5,
       rx_dout_reg_6,
       rx_dout_reg_7,
       rx_dout_reg_0,
       rx_dout_reg_1,
       rx_dout_reg_2,
       rx_byte_2,
       rx_byte_1,
       rx_byte_0,
       rx_byte_7,
       rx_byte_6,
       rx_byte_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreUARTapb_2_0_OVERFLOW,
       CoreUARTapb_2_0_RXRDY,
       N_669,
       N_432,
       CoreUARTapb_2_0_PARITY_ERR,
       CoreAPB3_0_APBmslave0_PENABLE,
       CoreAPB3_0_APBmslave0_PWRITE,
       clear_overflow_0_a2_0_0,
       N_423,
       N_367,
       mss_sb_0_TX,
       CoreUARTapb_2_0_TXRDY,
       Echo_control_0_TX,
       CoreUARTapb_2_0_FRAMING_ERR
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [4:3] data_out;
input  [2:2] CoreAPB3_0_APBmslave0_PADDR;
input  [7:0] controlReg1;
input  [7:0] controlReg2;
output rx_dout_reg_5;
output rx_dout_reg_6;
output rx_dout_reg_7;
output rx_dout_reg_0;
output rx_dout_reg_1;
output rx_dout_reg_2;
output rx_byte_2;
output rx_byte_1;
output rx_byte_0;
output rx_byte_7;
output rx_byte_6;
output rx_byte_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output CoreUARTapb_2_0_OVERFLOW;
output CoreUARTapb_2_0_RXRDY;
output N_669;
input  N_432;
output CoreUARTapb_2_0_PARITY_ERR;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  CoreAPB3_0_APBmslave0_PWRITE;
output clear_overflow_0_a2_0_0;
input  N_423;
input  N_367;
output mss_sb_0_TX;
output CoreUARTapb_2_0_TXRDY;
input  Echo_control_0_TX;
output CoreUARTapb_2_0_FRAMING_ERR;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, 
        \rx_dout_reg[3]_net_1 , VCC_net_1, \rx_dout[3] , 
        rx_dout_reg4_i_0, GND_net_1, \rx_dout_reg[4]_net_1 , 
        \rx_dout[4] , \rx_dout[5] , \rx_dout[6] , \rx_dout[7] , 
        \tx_hold_reg[0]_net_1 , tx_hold_reg5, \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[4]_net_1 , \tx_hold_reg[5]_net_1 , 
        \tx_hold_reg[6]_net_1 , \tx_hold_reg[7]_net_1 , \rx_dout[0] , 
        \rx_dout[1] , \rx_dout[2] , \rx_state[0]_net_1 , 
        \rx_state_ns[0] , \rx_state[1]_net_1 , N_91_i, rx_dout_reg4, 
        rx_dout_reg_empty_1_sqmuxa_i_0, overflow_reg5, 
        un1_clear_overflow_0_net_1, RXRDY5, clear_parity_reg_net_1, 
        clear_parity_reg0, clear_parity_en, fifo_write_tx_net_1, 
        tx_hold_reg5_i_0, fifo_full_rx, fifo_write, N_347_i_0, 
        \rx_byte_in[2] , \rx_byte_in[1] , \rx_byte_in[0] , 
        \rx_byte[4] , \rx_byte_in[4]_net_1 , \rx_byte_in[7]_net_1 , 
        \rx_byte_in[6]_net_1 , \rx_byte_in[5]_net_1 , \rx_byte[3] , 
        \rx_byte_in[3]_net_1 , rx_idle, stop_strobe, 
        fifo_write_rx_1_i_a2_0_a2_net_1, fifo_empty_rx, xmit_clock, 
        baud_clock, N_289, \tx_dout_reg[0] , \tx_dout_reg[1] , 
        \tx_dout_reg[2] , \tx_dout_reg[3] , \tx_dout_reg[4] , 
        \tx_dout_reg[5] , \tx_dout_reg[6] , \tx_dout_reg[7] , 
        fifo_read_tx, fifo_read_tx_i_0, fifo_full_tx_i_0, 
        fifo_empty_tx;
    
    SLE \tx_hold_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[5]_net_1 ));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_0));
    CFG3 #( .INIT(8'h01) )  fifo_write_rx_1_i_a2_0_a2 (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(fifo_write_rx_1_i_a2_0_a2_net_1));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2_0[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    mss_sb_CoreUARTapb_2_0_Rx_async_1s_0s_1s_2s make_RX (.rx_byte({
        rx_byte_7, rx_byte_6, rx_byte_5, \rx_byte[4] , \rx_byte[3] , 
        rx_byte_2, rx_byte_1, rx_byte_0}), .controlReg2({
        controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .clear_parity_reg(clear_parity_reg_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), 
        .Echo_control_0_TX(Echo_control_0_TX), 
        .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR), 
        .stop_strobe(stop_strobe), .CoreUARTapb_2_0_FRAMING_ERR(
        CoreUARTapb_2_0_FRAMING_ERR), .clear_parity_en(clear_parity_en)
        , .fifo_write(fifo_write), .rx_idle(rx_idle));
    SLE \tx_hold_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[0]_net_1 ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[3]_net_1 ));
    mss_sb_CoreUARTapb_2_0_fifo_256x8 \genblk2.tx_fifo  (.tx_dout_reg({
        \tx_dout_reg[7] , \tx_dout_reg[6] , \tx_dout_reg[5] , 
        \tx_dout_reg[4] , \tx_dout_reg[3] , \tx_dout_reg[2] , 
        \tx_dout_reg[1] , \tx_dout_reg[0] }), .tx_hold_reg({
        \tx_hold_reg[7]_net_1 , \tx_hold_reg[6]_net_1 , 
        \tx_hold_reg[5]_net_1 , \tx_hold_reg[4]_net_1 , 
        \tx_hold_reg[3]_net_1 , \tx_hold_reg[2]_net_1 , 
        \tx_hold_reg[1]_net_1 , \tx_hold_reg[0]_net_1 }), 
        .fifo_write_tx(fifo_write_tx_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[3]  (.A(\rx_byte[3] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[3]_net_1 ), .Y(
        data_out[3]));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE clear_framing_error_reg0 (.D(clear_parity_en), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(clear_parity_reg0));
    SLE \tx_hold_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3_0_x2[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_91_i));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(GL0_INST), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[5]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_5), .Y(
        \rx_byte_in[5]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in_0_a2[0]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_0), .Y(\rx_byte_in[0] )
        );
    CFG4 #( .INIT(16'h4000) )  \reg_write.tx_hold_reg5_0_a2_0  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .C(
        CoreAPB3_0_APBmslave0_PENABLE), .D(N_423), .Y(N_669));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[4]  (.A(\rx_byte[4] ), .B(
        CoreUARTapb_2_0_PARITY_ERR), .C(\rx_dout_reg[4]_net_1 ), .Y(
        data_out[4]));
    mss_sb_CoreUARTapb_2_0_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s make_TX (
        .tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .controlReg2({controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .N_289(N_289)
        , .mss_sb_0_TX(mss_sb_0_TX), .CoreUARTapb_2_0_TXRDY(
        CoreUARTapb_2_0_TXRDY), .fifo_full_tx_i_0(fifo_full_tx_i_0), 
        .xmit_clock(xmit_clock), .baud_clock(baud_clock), 
        .fifo_empty_tx(fifo_empty_tx));
    CFG3 #( .INIT(8'hFE) )  \genblk1.RXRDY5_0  (.A(rx_idle), .B(
        stop_strobe), .C(rx_dout_reg_empty_net_1), .Y(RXRDY5));
    SLE \tx_hold_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[6]_net_1 ));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \reg_write.tx_hold_reg5_0_a2  (.A(N_669), 
        .B(N_432), .Y(tx_hold_reg5));
    mss_sb_CoreUARTapb_2_0_Clock_gen_0s make_CLOCK_GEN (.controlReg1({
        controlReg1[7], controlReg1[6], controlReg1[5], controlReg1[4], 
        controlReg1[3], controlReg1[2], controlReg1[1], controlReg1[0]})
        , .controlReg2({controlReg2[7], controlReg2[6], controlReg2[5], 
        controlReg2[4], controlReg2[3]}), .xmit_clock(xmit_clock), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .N_289(N_289));
    SLE \rx_state[1]  (.D(N_91_i), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_7));
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_1));
    SLE clear_parity_reg (.D(clear_parity_reg0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_reg_net_1));
    CFG2 #( .INIT(4'h7) )  \reg_write.tx_hold_reg5_0_a2_i  (.A(N_669), 
        .B(N_432), .Y(tx_hold_reg5_i_0));
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_5));
    SLE overflow_reg (.D(overflow_reg5), .CLK(GL0_INST), .EN(
        un1_clear_overflow_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_0_OVERFLOW));
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_6));
    CFG2 #( .INIT(4'h2) )  clear_overflow_0_a2_0_0_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PENABLE), .B(
        CoreAPB3_0_APBmslave0_PWRITE), .Y(clear_overflow_0_a2_0_0));
    CFG4 #( .INIT(16'hECCC) )  un1_clear_overflow_0 (.A(
        clear_overflow_0_a2_0_0), .B(overflow_reg5), .C(N_432), .D(
        N_367), .Y(un1_clear_overflow_0_net_1));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \tx_hold_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[7]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(GL0_INST), 
        .EN(RXRDY5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_0_RXRDY));
    mss_sb_CoreUARTapb_2_0_fifo_256x8_0 \genblk3.rx_fifo  (.rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_state({\rx_state[1]_net_1 , \rx_state[0]_net_1 }), 
        .rx_byte_in({\rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte_in[4]_net_1 , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[2] , \rx_byte_in[1] , 
        \rx_byte_in[0] }), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .fifo_write_rx_1_i_a2_0_a2(fifo_write_rx_1_i_a2_0_a2_net_1), 
        .N_347_i_0(N_347_i_0), .rx_dout_reg_empty(
        rx_dout_reg_empty_net_1), .fifo_empty_rx(fifo_empty_rx), 
        .fifo_full_rx(fifo_full_rx));
    SLE \tx_hold_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in_0_a2[2]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_2), .Y(\rx_byte_in[2] )
        );
    CFG2 #( .INIT(4'h4) )  \rx_byte_in_0_a2[1]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_1), .Y(\rx_byte_in[1] )
        );
    SLE fifo_write_tx (.D(tx_hold_reg5_i_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_write_tx_net_1));
    CFG3 #( .INIT(8'hFE) )  fifo_write_rx_1_i_a2_0_a2_i (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(N_347_i_0));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[6]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_6), .Y(
        \rx_byte_in[6]_net_1 ));
    CFG2 #( .INIT(4'h2) )  overflow_reg5_0_a2_0_a2 (.A(fifo_full_rx), 
        .B(fifo_write), .Y(overflow_reg5));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[7]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(rx_byte_7), .Y(
        \rx_byte_in[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[3]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[3] ), .Y(
        \rx_byte_in[3]_net_1 ));
    SLE \tx_hold_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hB333) )  rx_dout_reg_empty_1_sqmuxa_i (.A(
        clear_overflow_0_a2_0_0), .B(rx_dout_reg4), .C(N_432), .D(
        N_367), .Y(rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_2));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[4]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(\rx_byte[4] ), .Y(
        \rx_byte_in[4]_net_1 ));
    SLE \tx_hold_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[4]_net_1 ));
    
endmodule


module 
        mss_sb_CoreUARTapb_2_0_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s(
        
       CoreAPB3_0_APBmslave0_PWDATA,
       CoreAPB3_0_APBmslave2_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_423,
       N_99_1,
       N_367,
       CoreUARTapb_2_0_PARITY_ERR,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE,
       psh_negedge_reg_1_sqmuxa_6_2,
       N_432,
       N_437,
       CoreUARTapb_2_0_RXRDY,
       CoreUARTapb_2_0_TXRDY,
       CoreUARTapb_2_0_FRAMING_ERR,
       CoreUARTapb_2_0_OVERFLOW,
       N_669,
       clear_overflow_0_a2_0_0,
       mss_sb_0_TX,
       Echo_control_0_TX
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [7:0] CoreAPB3_0_APBmslave2_PRDATA;
input  [4:2] CoreAPB3_0_APBmslave0_PADDR;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output N_423;
output N_99_1;
output N_367;
output CoreUARTapb_2_0_PARITY_ERR;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  psh_negedge_reg_1_sqmuxa_6_2;
input  N_432;
input  N_437;
output CoreUARTapb_2_0_RXRDY;
output CoreUARTapb_2_0_TXRDY;
output CoreUARTapb_2_0_FRAMING_ERR;
output CoreUARTapb_2_0_OVERFLOW;
output N_669;
output clear_overflow_0_a2_0_0;
output mss_sb_0_TX;
input  Echo_control_0_TX;

    wire \controlReg1[4]_net_1 , VCC_net_1, controlReg14, GND_net_1, 
        \controlReg1[5]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[7]_net_1 , \NxtPrdata[5] , N_422, \NxtPrdata[6] , 
        \NxtPrdata[7] , \controlReg2[0]_net_1 , controlReg24, 
        \controlReg2[1]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[7]_net_1 , \controlReg1[0]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[3]_net_1 , \NxtPrdata[0] , \NxtPrdata[1] , 
        \NxtPrdata[2] , \NxtPrdata[3] , \NxtPrdata[4] , 
        \NxtPrdata_5_bm_0[3] , \NxtPrdata_5_am_0[3] , 
        \NxtPrdata_5_bm_1[4] , \NxtPrdata_5_am_1[4] , 
        \NxtPrdata_5_bm_1[7] , \NxtPrdata_5_am_1[7] , 
        \NxtPrdata_5_bm_1[5] , \NxtPrdata_5_am_1[5] , 
        \NxtPrdata_5_bm_0[6] , \NxtPrdata_5_am_0[6] , N_153, N_344, 
        N_341, N_338, \rx_byte[0] , \rx_dout_reg[0] , N_345, 
        \rx_byte[1] , \rx_dout_reg[1] , N_342, \rx_byte[2] , 
        \rx_dout_reg[2] , N_339, \rx_dout_reg[6] , \rx_byte[6] , 
        \rx_dout_reg[5] , \rx_byte[5] , \rx_dout_reg[7] , \rx_byte[7] , 
        \data_out[4] , \data_out[3] ;
    
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[4]  (.A(
        CoreUARTapb_2_0_FRAMING_ERR), .B(\data_out[4] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_1[4] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[5]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[5] ), 
        .D(\rx_byte[5] ), .Y(\NxtPrdata_5_am_1[5] ));
    SLE \controlReg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[5]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \NxtPrdata_5_0[0]  (.A(
        CoreUARTapb_2_0_TXRDY), .B(N_153), .C(N_344), .D(N_345), .Y(
        \NxtPrdata[0] ));
    SLE \controlReg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[7]_net_1 ));
    SLE \iPRDATA[1]  (.D(\NxtPrdata[1] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[1]));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[6]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[6] ), 
        .D(\rx_byte[6] ), .Y(\NxtPrdata_5_am_0[6] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[7]  (.A(
        \controlReg2[7]_net_1 ), .B(\controlReg1[7]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_1[7] ));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[1]  (.A(
        \controlReg1[1]_net_1 ), .B(\controlReg2[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_341));
    SLE \controlReg2[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[4]_net_1 ));
    SLE \iPRDATA[4]  (.D(\NxtPrdata[4] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[4]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_0[2]  (.A(
        \rx_byte[2] ), .B(\rx_dout_reg[2] ), .C(N_367), .D(
        CoreUARTapb_2_0_PARITY_ERR), .Y(N_339));
    SLE \iPRDATA[3]  (.D(\NxtPrdata[3] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[3]));
    SLE \controlReg2[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[6]_net_1 ));
    SLE \controlReg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[4]  (.A(
        \controlReg2[4]_net_1 ), .B(\controlReg1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_1[4] ));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_0[0]  (.A(
        \rx_byte[0] ), .B(\rx_dout_reg[0] ), .C(N_367), .D(
        CoreUARTapb_2_0_PARITY_ERR), .Y(N_345));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[3]  (.A(
        CoreUARTapb_2_0_OVERFLOW), .B(\data_out[3] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[3] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[5]  (.A(
        \controlReg2[5]_net_1 ), .B(\controlReg1[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_1[5] ));
    CFG2 #( .INIT(4'h2) )  \NxtPrdata_3_1[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_99_1));
    SLE \controlReg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[6]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \NxtPrdata_5_0_a2_4[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_423));
    SLE \controlReg2[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[3]_net_1 ));
    SLE \controlReg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[2]_net_1 ));
    SLE \controlReg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[4]_net_1 ));
    SLE \iPRDATA[5]  (.D(\NxtPrdata[5] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[5]));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[0]  (.A(
        \controlReg1[0]_net_1 ), .B(\controlReg2[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_344));
    SLE \iPRDATA[7]  (.D(\NxtPrdata[7] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[7]));
    SLE \controlReg2[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24_0_a2  (.A(
        N_432), .B(CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(
        controlReg24));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[6]  (.A(
        \controlReg2[6]_net_1 ), .B(\controlReg1[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[6] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_1[4] ), .C(
        \NxtPrdata_5_am_1[4] ), .Y(\NxtPrdata[4] ));
    SLE \controlReg2[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[7]_net_1 ));
    SLE \iPRDATA[2]  (.D(\NxtPrdata[2] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[2]));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[3] ), .C(
        \NxtPrdata_5_am_0[3] ), .Y(\NxtPrdata[3] ));
    SLE \controlReg2[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[5]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[3]  (.A(
        \controlReg2[3]_net_1 ), .B(\controlReg1[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[3] ));
    SLE \controlReg2[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[2]_net_1 ));
    CFG4 #( .INIT(16'hA0C0) )  \NxtPrdata_5_0_a2_0[1]  (.A(
        \rx_byte[1] ), .B(\rx_dout_reg[1] ), .C(N_367), .D(
        CoreUARTapb_2_0_PARITY_ERR), .Y(N_342));
    SLE \iPRDATA[6]  (.D(\NxtPrdata[6] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[6]));
    SLE \iPRDATA[0]  (.D(\NxtPrdata[0] ), .CLK(GL0_INST), .EN(N_422), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PRDATA[0]));
    mss_sb_CoreUARTapb_2_0_COREUART_1s_1s_0s_15s_0s uUART (
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .data_out({\data_out[4] , 
        \data_out[3] }), .CoreAPB3_0_APBmslave0_PADDR({
        CoreAPB3_0_APBmslave0_PADDR[2]}), .controlReg1({
        \controlReg1[7]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[5]_net_1 , \controlReg1[4]_net_1 , 
        \controlReg1[3]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[0]_net_1 }), .controlReg2({
        \controlReg2[7]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[1]_net_1 , \controlReg2[0]_net_1 }), 
        .rx_dout_reg_5(\rx_dout_reg[5] ), .rx_dout_reg_6(
        \rx_dout_reg[6] ), .rx_dout_reg_7(\rx_dout_reg[7] ), 
        .rx_dout_reg_0(\rx_dout_reg[0] ), .rx_dout_reg_1(
        \rx_dout_reg[1] ), .rx_dout_reg_2(\rx_dout_reg[2] ), 
        .rx_byte_2(\rx_byte[2] ), .rx_byte_1(\rx_byte[1] ), .rx_byte_0(
        \rx_byte[0] ), .rx_byte_7(\rx_byte[7] ), .rx_byte_6(
        \rx_byte[6] ), .rx_byte_5(\rx_byte[5] ), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .CoreUARTapb_2_0_OVERFLOW(
        CoreUARTapb_2_0_OVERFLOW), .CoreUARTapb_2_0_RXRDY(
        CoreUARTapb_2_0_RXRDY), .N_669(N_669), .N_432(N_432), 
        .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .clear_overflow_0_a2_0_0(clear_overflow_0_a2_0_0), .N_423(
        N_423), .N_367(N_367), .mss_sb_0_TX(mss_sb_0_TX), 
        .CoreUARTapb_2_0_TXRDY(CoreUARTapb_2_0_TXRDY), 
        .Echo_control_0_TX(Echo_control_0_TX), 
        .CoreUARTapb_2_0_FRAMING_ERR(CoreUARTapb_2_0_FRAMING_ERR));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_1[7] ), .C(
        \NxtPrdata_5_am_1[7] ), .Y(\NxtPrdata[7] ));
    CFG4 #( .INIT(16'hCA00) )  \NxtPrdata_5_0_a2[2]  (.A(
        \controlReg1[2]_net_1 ), .B(\controlReg2[2]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_338));
    CFG4 #( .INIT(16'hFFF8) )  \NxtPrdata_5_0[2]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_153), .C(N_338), .D(N_339), 
        .Y(\NxtPrdata[2] ));
    CFG3 #( .INIT(8'h04) )  \NxtPrdata_5_0_a2_3[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_153));
    CFG3 #( .INIT(8'h10) )  \NxtPrdata_5_0_a2_2[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_367));
    SLE \controlReg2[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[0]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[6] ), .C(
        \NxtPrdata_5_am_0[6] ), .Y(\NxtPrdata[6] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[7]  (.A(
        CoreUARTapb_2_0_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[7] ), 
        .D(\rx_byte[7] ), .Y(\NxtPrdata_5_am_1[7] ));
    SLE \controlReg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[1]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \p_CtrlReg1Seq.controlReg14_0_a2  (.A(
        N_432), .B(CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(
        controlReg14));
    CFG4 #( .INIT(16'h0100) )  un1_NxtPrdata23_i_a2 (.A(
        CoreAPB3_0_APBmslave0_PWRITE), .B(
        CoreAPB3_0_APBmslave0_PENABLE), .C(
        psh_negedge_reg_1_sqmuxa_6_2), .D(N_432), .Y(N_422));
    CFG4 #( .INIT(16'hFFF8) )  \NxtPrdata_5_0[1]  (.A(
        CoreUARTapb_2_0_RXRDY), .B(N_153), .C(N_341), .D(N_342), .Y(
        \NxtPrdata[1] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_1[5] ), .C(
        \NxtPrdata_5_am_1[5] ), .Y(\NxtPrdata[5] ));
    SLE \controlReg1[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[0]_net_1 ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Rx_async_1s_0s_1s_2s(
       rx_byte,
       rx_state,
       controlReg2,
       clear_parity_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       GPS_TX_c,
       CoreUARTapb_2_1_PARITY_ERR,
       stop_strobe,
       CoreUARTapb_2_1_FRAMING_ERR,
       clear_parity_en,
       fifo_write
    );
output [7:0] rx_byte;
output [1:0] rx_state;
input  [2:0] controlReg2;
input  clear_parity_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  baud_clock;
input  GPS_TX_c;
output CoreUARTapb_2_1_PARITY_ERR;
output stop_strobe;
output CoreUARTapb_2_1_FRAMING_ERR;
output clear_parity_en;
output fifo_write;

    wire clear_parity_reg_i_0, \rx_bit_cnt[0]_net_1 , VCC_net_1, 
        \rx_bit_cnt_4[0] , GND_net_1, \rx_bit_cnt[1]_net_1 , 
        \rx_bit_cnt_4[1] , \rx_bit_cnt[2]_net_1 , \rx_bit_cnt_4[2] , 
        \rx_bit_cnt[3]_net_1 , \rx_bit_cnt_4[3] , \samples[1]_net_1 , 
        \samples[2]_net_1 , \rx_shift[0]_net_1 , \rx_shift_11[0] , 
        un1_samples7_1_0_1, \rx_shift[1]_net_1 , \rx_shift_11[1] , 
        \rx_shift[2]_net_1 , \rx_shift_11[2] , \rx_shift[3]_net_1 , 
        \rx_shift_11[3] , \rx_shift[4]_net_1 , \rx_shift_11[4] , 
        \rx_shift[5]_net_1 , \rx_shift_11[5] , \rx_shift[6]_net_1 , 
        \rx_shift_11[6] , \rx_shift[7]_net_1 , \rx_shift_11[7] , 
        \rx_shift[8]_net_1 , \rx_shift_11[8] , 
        \receive_count[0]_net_1 , \receive_count_3[0] , 
        \receive_count[1]_net_1 , \receive_count_3[1] , 
        \receive_count[2]_net_1 , \receive_count_3[2] , 
        \receive_count[3]_net_1 , \receive_count_3[3] , 
        clear_parity_en_9, \rx_byte_2[7] , \samples[0]_net_1 , N_310, 
        parity_err_1_sqmuxa_i_0, rx_parity_calc_net_1, 
        rx_parity_calc_4, framing_error_int_net_1, 
        framing_error_int_0_sqmuxa_net_1, N_238, 
        framing_error_1_sqmuxa_i_0, N_233_i_0, \rx_state_ns[0] , 
        clear_parity_en_9_i_0, framing_error_int10, CO1, 
        rx_bit_cnt_0_sqmuxa, rx_state19_li, 
        un1_parity_err_0_sqmuxa_2_1_0_net_1, 
        un1_parity_err_0_sqmuxa_2_1_net_1, un1_parity_err31_0_net_1, 
        N_238_1, N_242, framing_error_int_0_sqmuxa_1_net_1, rx_state10, 
        rx_state19_0, framing_error_int5, rx_state19_NE_1, 
        rx_parity_calc4, rx_bit_cnt_1_sqmuxa, \rx_shift_9[8] , 
        \rx_shift_9[7] , \rx_shift_9[6] , receive_count8;
    
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  framing_error_int_2_sqmuxa_0_a3 (.A(
        framing_error_int10), .B(rx_state[1]), .Y(N_238));
    CFG3 #( .INIT(8'hF8) )  un1_samples7_1_0 (.A(baud_clock), .B(
        framing_error_int10), .C(rx_bit_cnt_0_sqmuxa), .Y(
        un1_samples7_1_0_1));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[0]));
    CFG4 #( .INIT(16'h8000) )  framing_error_int_0_sqmuxa (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        framing_error_int5), .D(framing_error_int_0_sqmuxa_1_net_1), 
        .Y(framing_error_int_0_sqmuxa_net_1));
    SLE \receive_count[1]  (.D(\receive_count_3[1] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[1]_net_1 ));
    SLE \rx_shift[7]  (.D(\rx_shift_11[7] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \rx_par_calc.rx_parity_calc4  (.A(
        framing_error_int10), .B(controlReg2[1]), .Y(rx_parity_calc4));
    CFG4 #( .INIT(16'h1441) )  
        \make_parity_err.parity_err_12_iv_0_111_a2  (.A(
        clear_parity_reg), .B(framing_error_int5), .C(
        rx_parity_calc_net_1), .D(controlReg2[2]), .Y(N_310));
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[0]_net_1 ));
    CFG4 #( .INIT(16'h72F0) )  \receive_shift.rx_shift_11_RNO[8]  (.A(
        controlReg2[1]), .B(framing_error_int5), .C(
        \rx_shift[8]_net_1 ), .D(controlReg2[0]), .Y(\rx_shift_9[8] ));
    CFG3 #( .INIT(8'h40) )  
        \receive_full_indicator.clear_parity_en_9_0_a3  (.A(
        rx_state19_li), .B(rx_state[0]), .C(baud_clock), .Y(
        clear_parity_en_9));
    CFG2 #( .INIT(4'h1) )  \rcv_cnt.receive_count_3[0]  (.A(
        receive_count8), .B(\receive_count[0]_net_1 ), .Y(
        \receive_count_3[0] ));
    CFG1 #( .INIT(2'h1) )  framing_error_RNO (.A(clear_parity_reg), .Y(
        clear_parity_reg_i_0));
    CFG3 #( .INIT(8'h06) )  \rcv_cnt.receive_count_3[1]  (.A(
        \receive_count[1]_net_1 ), .B(\receive_count[0]_net_1 ), .C(
        receive_count8), .Y(\receive_count_3[1] ));
    CFG3 #( .INIT(8'h14) )  \rcv_cnt.receive_count_3[2]  (.A(
        receive_count8), .B(\receive_count[2]_net_1 ), .C(N_238_1), .Y(
        \receive_count_3[2] ));
    CFG3 #( .INIT(8'h04) )  rx_bit_cnt_0_sqmuxa_0_a3 (.A(rx_state[1]), 
        .B(baud_clock), .C(rx_state[0]), .Y(rx_bit_cnt_0_sqmuxa));
    CFG4 #( .INIT(16'h90F6) )  \receive_shift.rx_shift_9_u[7]  (.A(
        controlReg2[0]), .B(controlReg2[1]), .C(N_242), .D(
        framing_error_int5), .Y(\rx_shift_9[7] ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[0]  (.A(
        \rx_shift[1]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(\receive_count_3[3] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[4]));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[8]  (.A(
        rx_state[1]), .B(\rx_shift_9[8] ), .C(rx_state[0]), .Y(
        \rx_shift_11[8] ));
    SLE rx_parity_calc (.D(rx_parity_calc_4), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_parity_calc_net_1));
    SLE \rx_bit_cnt[2]  (.D(\rx_bit_cnt_4[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[2]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[3]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(CO1), .D(
        rx_bit_cnt_0_sqmuxa), .Y(\rx_bit_cnt_4[3] ));
    CFG4 #( .INIT(16'h0002) )  \rcv_cnt.rx_state10_0_a3  (.A(
        \receive_count[3]_net_1 ), .B(\receive_count[2]_net_1 ), .C(
        \receive_count[1]_net_1 ), .D(\receive_count[0]_net_1 ), .Y(
        rx_state10));
    SLE \rx_bit_cnt[1]  (.D(\rx_bit_cnt_4[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[1]_net_1 ));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[7]  (.A(
        rx_state[1]), .B(\rx_shift_9[7] ), .C(rx_state[0]), .Y(
        \rx_shift_11[7] ));
    CFG3 #( .INIT(8'hAC) )  \receive_shift.rx_shift_9_0[7]  (.A(
        \rx_shift[8]_net_1 ), .B(\rx_shift[7]_net_1 ), .C(
        controlReg2[1]), .Y(N_242));
    CFG4 #( .INIT(16'hFFBD) )  \rcv_sm.rx_state19_NE_1  (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        \rx_bit_cnt[2]_net_1 ), .D(rx_state19_0), .Y(rx_state19_NE_1));
    SLE stop_strobe_inst_1 (.D(N_238), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG4 #( .INIT(16'h0C2E) )  \rx_state_RNO[1]  (.A(rx_state[0]), .B(
        rx_state[1]), .C(framing_error_int10), .D(rx_state19_li), .Y(
        N_233_i_0));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[1]));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[2]  (.A(
        \rx_shift[3]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(\receive_count_3[2] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[2]_net_1 ));
    SLE clear_parity_en_1 (.D(clear_parity_en_9), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_en));
    CFG4 #( .INIT(16'h0180) )  un1_parity_err_0_sqmuxa_2_1 (.A(
        controlReg2[0]), .B(un1_parity_err_0_sqmuxa_2_1_0_net_1), .C(
        \rx_bit_cnt[3]_net_1 ), .D(\rx_bit_cnt[2]_net_1 ), .Y(
        un1_parity_err_0_sqmuxa_2_1_net_1));
    CFG4 #( .INIT(16'h8000) )  \un1_rx_bit_cnt_1.CO1  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        framing_error_int10), .D(baud_clock), .Y(CO1));
    SLE \rx_state[1]  (.D(N_233_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_state[1]));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[6]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h8000) )  \rx_state_ns_i_a3_0_3[1]  (.A(
        \receive_count[3]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[0]_net_1 ), .Y(
        framing_error_int10));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[4]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[3]  (.A(
        \rx_shift[4]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(\rx_byte_2[7] ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[7]));
    CFG4 #( .INIT(16'hCFDE) )  \rcv_sm.rx_state19_NE  (.A(
        controlReg2[1]), .B(rx_state19_NE_1), .C(\rx_bit_cnt[3]_net_1 )
        , .D(controlReg2[0]), .Y(rx_state19_li));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[2]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(CO1), .Y(
        \rx_bit_cnt_4[2] ));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[3]));
    CFG2 #( .INIT(4'h8) )  rx_bit_cnt_1_sqmuxa_0_a3 (.A(
        framing_error_int10), .B(baud_clock), .Y(rx_bit_cnt_1_sqmuxa));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[2]));
    CFG2 #( .INIT(4'h8) )  \rcv_sm.rx_byte_2[7]  (.A(controlReg2[0]), 
        .B(\rx_shift[7]_net_1 ), .Y(\rx_byte_2[7] ));
    CFG3 #( .INIT(8'h2B) )  un1_parity_err_0_sqmuxa_2_1_0 (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[0]_net_1 ), .C(
        \rx_bit_cnt[1]_net_1 ), .Y(un1_parity_err_0_sqmuxa_2_1_0_net_1)
        );
    SLE parity_err (.D(N_310), .CLK(GL0_INST), .EN(
        parity_err_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_1_PARITY_ERR));
    SLE \rx_shift[6]  (.D(\rx_shift_11[6] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[6]_net_1 ));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[1]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[4]  (.A(
        \rx_shift[5]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[3]_net_1 ));
    CFG3 #( .INIT(8'hC8) )  \receive_shift.rx_shift_11[6]  (.A(
        rx_state[1]), .B(\rx_shift_9[6] ), .C(rx_state[0]), .Y(
        \rx_shift_11[6] ));
    SLE framing_error_int (.D(framing_error_int_0_sqmuxa_net_1), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(framing_error_int_net_1));
    CFG3 #( .INIT(8'h69) )  \rcv_sm.rx_state19_0  (.A(controlReg2[1]), 
        .B(\rx_bit_cnt[0]_net_1 ), .C(controlReg2[0]), .Y(rx_state19_0)
        );
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_state[0]));
    CFG4 #( .INIT(16'h1101) )  \rcv_cnt.receive_count8  (.A(
        rx_state[0]), .B(rx_state[1]), .C(framing_error_int5), .D(
        rx_state10), .Y(receive_count8));
    SLE \samples[2]  (.D(GPS_TX_c), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    CFG4 #( .INIT(16'h060C) )  \rcv_cnt.receive_count_3[3]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        receive_count8), .D(N_238_1), .Y(\receive_count_3[3] ));
    SLE \receive_count[0]  (.D(\receive_count_3[0] ), .CLK(GL0_INST), 
        .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[5]));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[5]  (.A(
        \rx_shift[6]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[5] ));
    CFG3 #( .INIT(8'hBF) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_i  (.A(
        rx_state19_li), .B(rx_state[0]), .C(baud_clock), .Y(
        clear_parity_en_9_i_0));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[0]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(
        rx_bit_cnt_1_sqmuxa), .Y(\rx_bit_cnt_4[0] ));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[5]_net_1 ));
    CFG4 #( .INIT(16'hBA10) )  \rx_state_ns_0[0]  (.A(rx_state[0]), .B(
        rx_state[1]), .C(rx_state10), .D(rx_state19_li), .Y(
        \rx_state_ns[0] ));
    CFG2 #( .INIT(4'h7) )  un1_parity_err31_0 (.A(baud_clock), .B(
        controlReg2[1]), .Y(un1_parity_err31_0_net_1));
    SLE \rx_bit_cnt[0]  (.D(\rx_bit_cnt_4[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[0]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  framing_error_1_sqmuxa_i (.A(
        framing_error_int_net_1), .B(clear_parity_reg), .C(baud_clock), 
        .Y(framing_error_1_sqmuxa_i_0));
    SLE \rx_shift[8]  (.D(\rx_shift_11[8] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \rx_state_ns_i_a3_0_1[1]  (.A(
        \receive_count[0]_net_1 ), .B(\receive_count[1]_net_1 ), .Y(
        N_238_1));
    CFG3 #( .INIT(8'hA8) )  \receive_shift.rx_shift_11[1]  (.A(
        \rx_shift[2]_net_1 ), .B(rx_state[0]), .C(rx_state[1]), .Y(
        \rx_shift_11[1] ));
    CFG3 #( .INIT(8'h40) )  framing_error_int_0_sqmuxa_1 (.A(
        \receive_count[0]_net_1 ), .B(rx_state[1]), .C(
        \receive_count[1]_net_1 ), .Y(
        framing_error_int_0_sqmuxa_1_net_1));
    CFG3 #( .INIT(8'h17) )  \rx_filtered.m3  (.A(\samples[1]_net_1 ), 
        .B(\samples[0]_net_1 ), .C(\samples[2]_net_1 ), .Y(
        framing_error_int5));
    SLE framing_error (.D(clear_parity_reg_i_0), .CLK(GL0_INST), .EN(
        framing_error_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_1_FRAMING_ERR));
    CFG4 #( .INIT(16'hF0B1) )  \receive_shift.rx_shift_11_RNO[6]  (.A(
        controlReg2[1]), .B(framing_error_int5), .C(
        \rx_shift[7]_net_1 ), .D(controlReg2[0]), .Y(\rx_shift_9[6] ));
    CFG4 #( .INIT(16'hAEAA) )  parity_err_1_sqmuxa_i (.A(
        clear_parity_reg), .B(framing_error_int10), .C(
        un1_parity_err31_0_net_1), .D(
        un1_parity_err_0_sqmuxa_2_1_net_1), .Y(parity_err_1_sqmuxa_i_0)
        );
    CFG4 #( .INIT(16'h2122) )  \rx_par_calc.rx_parity_calc_4_u  (.A(
        rx_parity_calc_net_1), .B(rx_state[1]), .C(framing_error_int5), 
        .D(rx_parity_calc4), .Y(rx_parity_calc_4));
    SLE \rx_bit_cnt[3]  (.D(\rx_bit_cnt_4[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[1]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        rx_bit_cnt_1_sqmuxa), .D(rx_bit_cnt_0_sqmuxa), .Y(
        \rx_bit_cnt_4[1] ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] tx_hold_reg;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), .C_WEN(
        INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), 
        .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_ctrl_128(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_3670_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, \counter[0]_net_1 , 
        VCC_net_1, un1_counter_cry_0_Y_4, GND_net_1, 
        \counter[1]_net_1 , un1_counter_cry_1_0_S_3, 
        \counter[2]_net_1 , un1_counter_cry_2_0_S_3, 
        \counter[3]_net_1 , un1_counter_cry_3_0_S_3, 
        \counter[4]_net_1 , un1_counter_cry_4_0_S_3, 
        \counter[5]_net_1 , un1_counter_cry_5_0_S_3, 
        \counter[6]_net_1 , un1_counter_s_6_S_3, \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \data_out_0[0] , 
        \data_out_0[1] , \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_308_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_309_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        empty_4_net_1, full_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_309_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_2_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[2]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S_3), .Y(), .FCO(
        un1_counter_cry_2));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_308 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_308_FCO));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_4_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[4]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S_3), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_308_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_3670_i_0 (.A(fifo_write_tx), .Y(
        N_3670_i_0_net_1));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[0]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  full_4_RNILIET (.A(\counter[0]_net_1 ), 
        .B(full_4_net_1), .C(\counter[6]_net_1 ), .D(
        \counter[5]_net_1 ), .Y(fifo_full_tx_i_0));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[6]));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_3_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[3]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S_3), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_309 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_309_FCO));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_tx), .C(fifo_write_tx), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_4), 
        .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_empty_tx));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNII4ID (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_3670_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_1_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_3), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_5_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[5]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S_3), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_1_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg({
        tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], 
        tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]})
        , .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_tx(fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(\counter[6]_net_1 ), 
        .FCI(un1_counter_cry_5), .S(un1_counter_s_6_S_3), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_256x8(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_1_fifo_ctrl_128 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.tx_dout_reg({
        tx_dout_reg[7], tx_dout_reg[6], tx_dout_reg[5], tx_dout_reg[4], 
        tx_dout_reg[3], tx_dout_reg[2], tx_dout_reg[1], tx_dout_reg[0]})
        , .tx_hold_reg({tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], 
        tx_hold_reg[4], tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], 
        tx_hold_reg[0]}), .fifo_write_tx(fifo_write_tx), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       controlReg2,
       fifo_read_tx,
       fifo_read_tx_i_0,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       xmit_pulse,
       GPS_RX_c,
       CoreUARTapb_2_1_TXRDY,
       fifo_full_tx_i_0,
       xmit_clock,
       baud_clock,
       fifo_empty_tx
    );
input  [7:0] tx_dout_reg;
input  [2:0] controlReg2;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  xmit_pulse;
output GPS_RX_c;
output CoreUARTapb_2_1_TXRDY;
input  fifo_full_tx_i_0;
input  xmit_clock;
input  baud_clock;
input  fifo_empty_tx;

    wire \tx_byte[4]_net_1 , VCC_net_1, N_133_i_0, GND_net_1, 
        \tx_byte[5]_net_1 , \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_122_i_0, \xmit_bit_sel[2]_net_1 , 
        N_124_i_0, \xmit_bit_sel[3]_net_1 , N_126_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , \tx_byte[2]_net_1 , 
        \tx_byte[3]_net_1 , tx_parity_net_1, tx_parity_5, 
        un1_tx_parity_1_sqmuxa_0_net_1, tx_4_iv_i_0, N_144_i_0, 
        \xmit_state_ns_i_0[6] , \xmit_state[6]_net_1 , 
        \xmit_state_ns[6] , \xmit_state[0]_net_1 , 
        \xmit_state_ns[0]_net_1 , \xmit_state[1]_net_1 , 
        \xmit_state[2]_net_1 , \xmit_state_ns[2]_net_1 , 
        \xmit_state[3]_net_1 , N_112_i_0, \xmit_state[4]_net_1 , 
        \xmit_state_ns[4]_net_1 , \xmit_state[5]_net_1 , 
        \xmit_state_ns[5]_net_1 , N_174, tx_2_u_am_1_1, tx_2_u_am, 
        tx_2_u_bm_1_1, tx_2_u_bm, tx_2, N_129, N_128_i, tx_3_i_m, 
        N_172, N_154;
    
    SLE tx_parity (.D(tx_parity_5), .CLK(GL0_INST), .EN(
        un1_tx_parity_1_sqmuxa_0_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_parity_net_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_1_TXRDY));
    CFG4 #( .INIT(16'h2000) )  \xmit_state_ns_a3[5]  (.A(
        \xmit_state[3]_net_1 ), .B(controlReg2[1]), .C(xmit_pulse), .D(
        N_172), .Y(N_154));
    CFG2 #( .INIT(4'h6) )  \xmit_state_ns_i_x2[3]  (.A(controlReg2[0]), 
        .B(\xmit_bit_sel[0]_net_1 ), .Y(N_128_i));
    SLE \xmit_state[3]  (.D(N_112_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[3]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \xmit_cnt.xmit_bit_sel_3_i_o2[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        N_129));
    CFG4 #( .INIT(16'h0031) )  \xmit_sel.tx_4_iv_i  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(tx_2), 
        .D(tx_3_i_m), .Y(tx_4_iv_i_0));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[0]_net_1 ));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[4]_net_1 ));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[0]_net_1 ), .B(\xmit_bit_sel[1]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_122_i_0));
    CFG4 #( .INIT(16'h8000) )  un1_tx_parity_1_sqmuxa_0_a2 (.A(
        \xmit_state[3]_net_1 ), .B(xmit_clock), .C(baud_clock), .D(
        controlReg2[1]), .Y(N_174));
    CFG2 #( .INIT(4'h8) )  \xmit_state_RNIHFLK[2]  (.A(xmit_pulse), .B(
        \xmit_state[2]_net_1 ), .Y(N_133_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNI2248 (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[5]_net_1 ));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[5]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(tx_2_u_bm_1_1), 
        .D(\xmit_bit_sel[1]_net_1 ), .Y(tx_2_u_bm));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(
        xmit_pulse), .Y(\xmit_state_ns[2]_net_1 ));
    CFG4 #( .INIT(16'hDC50) )  \xmit_state_ns[4]  (.A(xmit_pulse), .B(
        N_172), .C(\xmit_state[4]_net_1 ), .D(N_174), .Y(
        \xmit_state_ns[4]_net_1 ));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_126_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[3]_net_1 ));
    SLE \xmit_bit_sel[2]  (.D(N_124_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \xmit_sel.tx_2_u_ns  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(tx_2_u_bm), .C(tx_2_u_am), .Y(
        tx_2));
    SLE tx (.D(tx_4_iv_i_0), .CLK(GL0_INST), .EN(N_144_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(GPS_RX_c));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[3]_net_1 ));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[7]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_state_RNICRA11[1]  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(
        xmit_pulse), .D(\xmit_state[6]_net_1 ), .Y(N_144_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_bm_1_1));
    CFG2 #( .INIT(4'hE) )  un1_tx_parity_1_sqmuxa_0 (.A(N_174), .B(
        \xmit_state[5]_net_1 ), .Y(un1_tx_parity_1_sqmuxa_0_net_1));
    CFG4 #( .INIT(16'hF7A0) )  \xmit_state_RNO[3]  (.A(xmit_pulse), .B(
        N_172), .C(\xmit_state[2]_net_1 ), .D(\xmit_state[3]_net_1 ), 
        .Y(N_112_i_0));
    CFG3 #( .INIT(8'h06) )  \xmit_par_calc.tx_parity_5  (.A(tx_2), .B(
        tx_parity_net_1), .C(\xmit_state[5]_net_1 ), .Y(tx_parity_5));
    CFG4 #( .INIT(16'h0040) )  \xmit_state_ns_i_a2[3]  (.A(
        \xmit_bit_sel[3]_net_1 ), .B(\xmit_bit_sel[2]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(N_128_i), .Y(N_172));
    CFG3 #( .INIT(8'h82) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_state[3]_net_1 ), .B(N_129), .C(\xmit_bit_sel[2]_net_1 ), 
        .Y(N_124_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_am_1_1));
    CFG4 #( .INIT(16'hFDEC) )  \xmit_state_ns[5]  (.A(xmit_pulse), .B(
        N_154), .C(\xmit_state[4]_net_1 ), .D(\xmit_state[5]_net_1 ), 
        .Y(\xmit_state_ns[5]_net_1 ));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[6]_net_1 ));
    CFG3 #( .INIT(8'h82) )  \xmit_sel.tx_4_iv_i_RNO  (.A(
        \xmit_state[4]_net_1 ), .B(controlReg2[2]), .C(tx_parity_net_1)
        , .Y(tx_3_i_m));
    SLE \xmit_bit_sel[1]  (.D(N_122_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[1]_net_1 ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[1]_net_1 ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(GL0_INST), 
        .EN(xmit_pulse), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[2]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(tx_2_u_am_1_1), 
        .D(\xmit_bit_sel[1]_net_1 ), .Y(tx_2_u_am));
    CFG2 #( .INIT(4'h4) )  fifo_read_en0_1_i_a3 (.A(fifo_empty_tx), .B(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[6] ));
    SLE fifo_read_en0 (.D(\xmit_state_ns_i_0[6] ), .CLK(GL0_INST), .EN(
        N_144_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns[0]  (.A(fifo_empty_tx), 
        .B(xmit_pulse), .C(\xmit_state[5]_net_1 ), .D(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[0]_net_1 ));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[1]_net_1 ));
    SLE \xmit_state[4]  (.D(\xmit_state_ns[4]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[4]_net_1 ));
    CFG4 #( .INIT(16'h82A0) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_state[3]_net_1 ), .B(N_129), .C(\xmit_bit_sel[3]_net_1 ), 
        .D(\xmit_bit_sel[2]_net_1 ), .Y(N_126_i_0));
    SLE \xmit_state[6]  (.D(\xmit_state_ns[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[6]_net_1 ));
    CFG2 #( .INIT(4'hB) )  fifo_read_en0_1_i_a3_i (.A(fifo_empty_tx), 
        .B(\xmit_state[0]_net_1 ), .Y(\xmit_state_ns_i_0[6] ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_Clock_gen_0s(
       controlReg1,
       controlReg2,
       xmit_clock,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       xmit_pulse
    );
input  [7:0] controlReg1;
input  [7:3] controlReg2;
output xmit_clock;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output baud_clock;
output xmit_pulse;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNIURC7_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[4] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIM2N85[9]  (.A(
        VCC_net_1), .B(controlReg2[4]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[9] ), .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] )
        , .Y(), .FCO(\baud_cntr_cry[9] ));
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[1] ));
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[3] ));
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[3]_net_1 ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI61172[3]  (.A(
        VCC_net_1), .B(controlReg1[3]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[3] ), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] )
        , .Y(), .FCO(\baud_cntr_cry[3] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIE7M64[7]  (.A(
        VCC_net_1), .B(controlReg1[7]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[7] ), .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] )
        , .Y(), .FCO(\baud_cntr_cry[7] ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[9] ));
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNIURC7_Y), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(baud_clock));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIK58R5[10]  (.A(
        VCC_net_1), .B(controlReg2[5]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[10] ), .FCI(\baud_cntr_cry[9] ), .S(
        \baud_cntr_s[10] ), .Y(), .FCO(\baud_cntr_cry[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI6GR63[5]  (.A(
        VCC_net_1), .B(controlReg1[5]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[5] ), .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] )
        , .Y(), .FCO(\baud_cntr_cry[5] ));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[7] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI1KMN4[8]  (.A(
        VCC_net_1), .B(controlReg2[3]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[8] ), .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] )
        , .Y(), .FCO(\baud_cntr_cry[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIEQ671[1]  (.A(
        VCC_net_1), .B(controlReg1[1]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[1] ), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] )
        , .Y(), .FCO(\baud_cntr_cry[1] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[5] ));
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIKAPD6[11]  (.A(
        VCC_net_1), .B(controlReg2[6]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[11] ), .FCI(\baud_cntr_cry[10] ), .S(
        \baud_cntr_s[11] ), .Y(), .FCO(\baud_cntr_cry[11] ));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNIURC7  (.A(baud_cntr8_8)
        , .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(baud_cntr8_7), .FCI(
        VCC_net_1), .S(), .Y(baud_cntr8_1_RNIURC7_Y), .FCO(
        baud_cntr_cry_cy));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[0] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[10] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIPS3N1[2]  (.A(
        VCC_net_1), .B(controlReg1[2]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[2] ), .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] )
        , .Y(), .FCO(\baud_cntr_cry[2] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[6] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI5Q9N[0]  (.A(
        VCC_net_1), .B(controlReg1[0]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[0] ), .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), 
        .Y(), .FCO(\baud_cntr_cry[0] ));
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        xmit_clock));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h44700) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(controlReg2[7]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[12] ), .FCI(\baud_cntr_cry[11] ), .S(
        \baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[1]_net_1 ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIL7UM2[4]  (.A(
        VCC_net_1), .B(controlReg1[4]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[4] ), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] )
        , .Y(), .FCO(\baud_cntr_cry[4] ));
    CFG2 #( .INIT(4'h8) )  xmit_pulse_inst_1 (.A(baud_clock), .B(
        xmit_clock), .Y(xmit_pulse));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIPQOM3[6]  (.A(
        VCC_net_1), .B(controlReg1[6]), .C(baud_cntr8_1_RNIURC7_Y), .D(
        \baud_cntr[6] ), .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] )
        , .Y(), .FCO(\baud_cntr_cry[6] ));
    
endmodule


module mss_sb_CoreUARTapb_2_1_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte_in,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_rx_1
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte_in;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_rx_1;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte_in[7], rx_byte_in[6], 
        rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], 
        rx_byte_in[1], rx_byte_in[0]}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_rx_1), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_ctrl_128_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_3686_i_0,
       N_3687_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_3686_i_0;
input  N_3687_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_empty_rx;
output fifo_full_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[1]_net_1 , VCC_net_1, 
        un1_counter_cry_1_0_S_4, GND_net_1, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_4, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S_4, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_4, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_4, \counter[6]_net_1 , 
        un1_counter_s_6_S_4, \counter[0]_net_1 , un1_counter_cry_0_Y_3, 
        \data_out_0[0] , \data_out_0[1] , \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \wr_pointer[1]_net_1 , 
        \wr_pointer_s[1] , \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_310_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_311_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_4_net_1, empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_311_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIHD74 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_2_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[2]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_1), 
        .S(un1_counter_cry_2_0_S_4), .Y(), .FCO(un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(N_3686_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_4_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[4]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_3), 
        .S(un1_counter_cry_4_0_S_4), .Y(), .FCO(un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_310_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_310 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_310_FCO));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_4), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_3_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[3]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_2), 
        .S(un1_counter_cry_3_0_S_4), .Y(), .FCO(un1_counter_cry_3));
    ARI1 #( .INIT(20'h56699) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(GND_net_1), .S(), .Y(
        un1_counter_cry_0_Y_3), .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_empty_rx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_3687_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_1_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_4), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_311 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_311_FCO));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[1]));
    CFG4 #( .INIT(16'h8000) )  full (.A(\counter[0]_net_1 ), .B(
        full_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_full_rx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_5_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[5]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_4), 
        .S(un1_counter_cry_5_0_S_4), .Y(), .FCO(un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_1_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte_in({
        rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], 
        rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_rx_1(fifo_write_rx_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(
        \counter[6]_net_1 ), .FCI(un1_counter_cry_5), .S(
        un1_counter_s_6_S_4), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_3), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_1_fifo_256x8_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_3686_i_0,
       N_3687_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_empty_rx,
       fifo_full_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_3686_i_0;
input  N_3687_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_empty_rx;
output fifo_full_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_1_fifo_ctrl_128_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_byte_in({rx_byte_in[7], 
        rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], 
        rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_3686_i_0(N_3686_i_0), .N_3687_i_0(
        N_3687_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1), .fifo_empty_rx(
        fifo_empty_rx), .fifo_full_rx(fifo_full_rx));
    
endmodule


module mss_sb_CoreUARTapb_2_1_COREUART_1s_1s_0s_15s_0s(
       CoreAPB3_0_APBmslave0_PWDATA,
       data_out,
       controlReg1,
       controlReg2,
       rx_dout_reg_5,
       rx_dout_reg_6,
       rx_dout_reg_7,
       rx_byte_7,
       rx_byte_6,
       rx_byte_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreUARTapb_2_1_OVERFLOW,
       CoreUARTapb_2_1_RXRDY,
       N_669,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreUARTapb_2_1_PARITY_ERR,
       N_367,
       clear_overflow_0_a2_0_0,
       GPS_RX_c,
       CoreUARTapb_2_1_TXRDY,
       GPS_TX_c,
       CoreUARTapb_2_1_FRAMING_ERR
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [4:0] data_out;
input  [7:0] controlReg1;
input  [7:0] controlReg2;
output rx_dout_reg_5;
output rx_dout_reg_6;
output rx_dout_reg_7;
output rx_byte_7;
output rx_byte_6;
output rx_byte_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output CoreUARTapb_2_1_OVERFLOW;
output CoreUARTapb_2_1_RXRDY;
input  N_669;
input  CoreAPB3_0_APBmslave3_PSELx;
output CoreUARTapb_2_1_PARITY_ERR;
input  N_367;
input  clear_overflow_0_a2_0_0;
output GPS_RX_c;
output CoreUARTapb_2_1_TXRDY;
input  GPS_TX_c;
output CoreUARTapb_2_1_FRAMING_ERR;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, 
        \rx_dout_reg[3]_net_1 , VCC_net_1, \rx_dout[3] , 
        rx_dout_reg4_i_0, GND_net_1, \rx_dout_reg[4]_net_1 , 
        \rx_dout[4] , \rx_dout[5] , \rx_dout[6] , \rx_dout[7] , 
        \tx_hold_reg[0]_net_1 , tx_hold_reg5, \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[4]_net_1 , \tx_hold_reg[5]_net_1 , 
        \tx_hold_reg[6]_net_1 , \tx_hold_reg[7]_net_1 , 
        \rx_dout_reg[0]_net_1 , \rx_dout[0] , \rx_dout_reg[1]_net_1 , 
        \rx_dout[1] , \rx_dout_reg[2]_net_1 , \rx_dout[2] , 
        \rx_state[0]_net_1 , \rx_state_ns[0] , \rx_state[1]_net_1 , 
        N_143_i, rx_dout_reg4, rx_dout_reg_empty_1_sqmuxa_i_0, 
        overflow_reg5_net_1, un1_clear_overflow_net_1, RXRDY5, 
        clear_parity_reg_net_1, clear_parity_reg0, clear_parity_en, 
        fifo_write_tx_net_1, tx_hold_reg5_i_0, fifo_empty_rx, 
        N_3686_i_0, fifo_full_rx, fifo_write, N_3687_i_0, \rx_byte[4] , 
        \rx_byte_in[4]_net_1 , \rx_byte_in[7]_net_1 , \rx_byte[1] , 
        \rx_byte_in[1]_net_1 , \rx_byte[3] , \rx_byte_in[3]_net_1 , 
        \rx_byte[0] , \rx_byte_in[0]_net_1 , \rx_byte[2] , 
        \rx_byte_in[2]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , stop_strobe, \rx_state_0[1] , 
        \rx_state_0[0] , fifo_write_rx_1_net_1, fifo_read_rx_0_sqmuxa, 
        xmit_clock, baud_clock, xmit_pulse, \tx_dout_reg[0] , 
        \tx_dout_reg[1] , \tx_dout_reg[2] , \tx_dout_reg[3] , 
        \tx_dout_reg[4] , \tx_dout_reg[5] , \tx_dout_reg[6] , 
        \tx_dout_reg[7] , fifo_read_tx, fifo_read_tx_i_0, 
        fifo_full_tx_i_0, fifo_empty_tx;
    
    SLE \tx_hold_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  overflow_reg5 (.A(fifo_full_rx), .B(
        fifo_write), .Y(overflow_reg5_net_1));
    CFG3 #( .INIT(8'h01) )  fifo_write_rx_1_i (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(N_3687_i_0));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[0]_net_1 ));
    CFG4 #( .INIT(16'hFFFB) )  fifo_read_rx_0_sqmuxa_0_a2_i (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(N_3686_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_143_i));
    CFG3 #( .INIT(8'hFE) )  fifo_write_rx_1 (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(fifo_write_rx_1_net_1));
    mss_sb_CoreUARTapb_2_1_Rx_async_1s_0s_1s_2s make_RX (.rx_byte({
        rx_byte_7, rx_byte_6, rx_byte_5, \rx_byte[4] , \rx_byte[3] , 
        \rx_byte[2] , \rx_byte[1] , \rx_byte[0] }), .rx_state({
        \rx_state_0[1] , \rx_state_0[0] }), .controlReg2({
        controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .clear_parity_reg(clear_parity_reg_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .GPS_TX_c(
        GPS_TX_c), .CoreUARTapb_2_1_PARITY_ERR(
        CoreUARTapb_2_1_PARITY_ERR), .stop_strobe(stop_strobe), 
        .CoreUARTapb_2_1_FRAMING_ERR(CoreUARTapb_2_1_FRAMING_ERR), 
        .clear_parity_en(clear_parity_en), .fifo_write(fifo_write));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[1]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[1] ), .Y(
        \rx_byte_in[1]_net_1 ));
    SLE \tx_hold_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[3]_net_1 ));
    mss_sb_CoreUARTapb_2_1_fifo_256x8 \genblk2.tx_fifo  (.tx_dout_reg({
        \tx_dout_reg[7] , \tx_dout_reg[6] , \tx_dout_reg[5] , 
        \tx_dout_reg[4] , \tx_dout_reg[3] , \tx_dout_reg[2] , 
        \tx_dout_reg[1] , \tx_dout_reg[0] }), .tx_hold_reg({
        \tx_hold_reg[7]_net_1 , \tx_hold_reg[6]_net_1 , 
        \tx_hold_reg[5]_net_1 , \tx_hold_reg[4]_net_1 , 
        \tx_hold_reg[3]_net_1 , \tx_hold_reg[2]_net_1 , 
        \tx_hold_reg[1]_net_1 , \tx_hold_reg[0]_net_1 }), 
        .fifo_write_tx(fifo_write_tx_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[3]  (.A(\rx_byte[3] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[3]_net_1 ), .Y(
        data_out[3]));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE clear_framing_error_reg0 (.D(clear_parity_en), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(clear_parity_reg0));
    SLE \tx_hold_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(GL0_INST), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[5]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_5), .Y(
        \rx_byte_in[5]_net_1 ));
    CFG4 #( .INIT(16'hEEEF) )  \genblk1.RXRDY5  (.A(
        rx_dout_reg_empty_net_1), .B(stop_strobe), .C(\rx_state_0[1] ), 
        .D(\rx_state_0[0] ), .Y(RXRDY5));
    CFG4 #( .INIT(16'h0004) )  fifo_read_rx_0_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(
        fifo_read_rx_0_sqmuxa));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[4]  (.A(\rx_byte[4] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[4]_net_1 ), .Y(
        data_out[4]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[2]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[2] ), .Y(
        \rx_byte_in[2]_net_1 ));
    mss_sb_CoreUARTapb_2_1_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s make_TX (
        .tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .controlReg2({controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .xmit_pulse(
        xmit_pulse), .GPS_RX_c(GPS_RX_c), .CoreUARTapb_2_1_TXRDY(
        CoreUARTapb_2_1_TXRDY), .fifo_full_tx_i_0(fifo_full_tx_i_0), 
        .xmit_clock(xmit_clock), .baud_clock(baud_clock), 
        .fifo_empty_tx(fifo_empty_tx));
    SLE \tx_hold_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[6]_net_1 ));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \reg_write.tx_hold_reg5_0_a2  (.A(N_669), 
        .B(CoreAPB3_0_APBmslave3_PSELx), .Y(tx_hold_reg5));
    mss_sb_CoreUARTapb_2_1_Clock_gen_0s make_CLOCK_GEN (.controlReg1({
        controlReg1[7], controlReg1[6], controlReg1[5], controlReg1[4], 
        controlReg1[3], controlReg1[2], controlReg1[1], controlReg1[0]})
        , .controlReg2({controlReg2[7], controlReg2[6], controlReg2[5], 
        controlReg2[4], controlReg2[3]}), .xmit_clock(xmit_clock), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .xmit_pulse(
        xmit_pulse));
    SLE \rx_state[1]  (.D(N_143_i), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_7));
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  un1_clear_overflow (.A(N_367), .B(
        CoreAPB3_0_APBmslave3_PSELx), .C(overflow_reg5_net_1), .D(
        clear_overflow_0_a2_0_0), .Y(un1_clear_overflow_net_1));
    SLE clear_parity_reg (.D(clear_parity_reg0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_reg_net_1));
    CFG2 #( .INIT(4'h7) )  \reg_write.tx_hold_reg5_0_a2_i  (.A(N_669), 
        .B(CoreAPB3_0_APBmslave3_PSELx), .Y(tx_hold_reg5_i_0));
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_5));
    SLE overflow_reg (.D(overflow_reg5_net_1), .CLK(GL0_INST), .EN(
        un1_clear_overflow_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_1_OVERFLOW));
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[0]  (.A(\rx_byte[0] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[0]_net_1 ), .Y(
        data_out[0]));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[2]  (.A(\rx_byte[2] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[2]_net_1 ), .Y(
        data_out[2]));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_6));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \tx_hold_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[7]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(GL0_INST), 
        .EN(RXRDY5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_1_RXRDY));
    mss_sb_CoreUARTapb_2_1_fifo_256x8_0 \genblk3.rx_fifo  (.rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_byte_in({\rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte_in[4]_net_1 , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[1]_net_1 , \rx_byte_in[0]_net_1 }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_3686_i_0(N_3686_i_0), .N_3687_i_0(
        N_3687_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1_net_1), .fifo_empty_rx(
        fifo_empty_rx), .fifo_full_rx(fifo_full_rx));
    SLE \tx_hold_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[3]_net_1 ));
    SLE fifo_write_tx (.D(tx_hold_reg5_i_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_write_tx_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[6]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_6), .Y(
        \rx_byte_in[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[1]  (.A(\rx_byte[1] ), .B(
        CoreUARTapb_2_1_PARITY_ERR), .C(\rx_dout_reg[1]_net_1 ), .Y(
        data_out[1]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[7]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(rx_byte_7), .Y(
        \rx_byte_in[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[3]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[3] ), .Y(
        \rx_byte_in[3]_net_1 ));
    SLE \tx_hold_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[1]_net_1 ));
    CFG4 #( .INIT(16'h8F0F) )  rx_dout_reg_empty_1_sqmuxa_i (.A(N_367), 
        .B(CoreAPB3_0_APBmslave3_PSELx), .C(rx_dout_reg4), .D(
        clear_overflow_0_a2_0_0), .Y(rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[4]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[4] ), .Y(
        \rx_byte_in[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[0]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\rx_byte[0] ), .Y(
        \rx_byte_in[0]_net_1 ));
    SLE \tx_hold_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[4]_net_1 ));
    
endmodule


module 
        mss_sb_CoreUARTapb_2_1_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s(
        
       CoreAPB3_0_APBmslave0_PWDATA,
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_425,
       CoreUARTapb_2_1_OVERFLOW,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE,
       psh_negedge_reg_1_sqmuxa_6_2,
       CoreAPB3_0_APBmslave3_PSELx,
       N_437,
       CoreUARTapb_2_1_PARITY_ERR,
       N_99_1,
       N_367,
       CoreUARTapb_2_1_FRAMING_ERR,
       CoreUARTapb_2_1_RXRDY,
       CoreUARTapb_2_1_TXRDY,
       N_669,
       clear_overflow_0_a2_0_0,
       GPS_RX_c,
       GPS_TX_c
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [4:2] CoreAPB3_0_APBmslave0_PADDR;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output N_425;
output CoreUARTapb_2_1_OVERFLOW;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;
input  psh_negedge_reg_1_sqmuxa_6_2;
input  CoreAPB3_0_APBmslave3_PSELx;
input  N_437;
output CoreUARTapb_2_1_PARITY_ERR;
input  N_99_1;
input  N_367;
output CoreUARTapb_2_1_FRAMING_ERR;
output CoreUARTapb_2_1_RXRDY;
output CoreUARTapb_2_1_TXRDY;
input  N_669;
input  clear_overflow_0_a2_0_0;
output GPS_RX_c;
input  GPS_TX_c;

    wire \controlReg1[4]_net_1 , VCC_net_1, controlReg14, GND_net_1, 
        \controlReg1[5]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[7]_net_1 , \NxtPrdata[5] , 
        un1_NxtPrdata23_i_a2_net_1, \NxtPrdata[6] , \NxtPrdata[7] , 
        \controlReg2[0]_net_1 , controlReg24, \controlReg2[1]_net_1 , 
        \controlReg2[2]_net_1 , \controlReg2[3]_net_1 , 
        \controlReg2[4]_net_1 , \controlReg2[5]_net_1 , 
        \controlReg2[6]_net_1 , \controlReg2[7]_net_1 , 
        \controlReg1[0]_net_1 , \controlReg1[1]_net_1 , 
        \controlReg1[2]_net_1 , \controlReg1[3]_net_1 , \NxtPrdata[0] , 
        \NxtPrdata[1] , \NxtPrdata[2] , \NxtPrdata[3] , \NxtPrdata[4] , 
        \NxtPrdata_5_bm[2]_net_1 , \NxtPrdata_5_am[2]_net_1 , 
        \NxtPrdata_5_bm_0[0] , \NxtPrdata_5_am_0[0] , 
        \NxtPrdata_5_bm[1]_net_1 , \NxtPrdata_5_am[1]_net_1 , 
        \NxtPrdata_5_bm_0[4] , \NxtPrdata_5_am_0[4] , 
        \NxtPrdata_5_bm_0[5] , \NxtPrdata_5_am_0[5] , 
        \NxtPrdata_5_bm_1[6] , \NxtPrdata_5_am_1[6] , 
        \NxtPrdata_5_bm_0[7] , \NxtPrdata_5_am_0[7] , N_608, N_606, 
        \rx_dout_reg[7] , \rx_byte[7] , \rx_dout_reg[6] , \rx_byte[6] , 
        \rx_dout_reg[5] , \rx_byte[5] , \data_out[3] , \data_out[4] , 
        \data_out[1] , \data_out[0] , \data_out[2] ;
    
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[4]  (.A(
        CoreUARTapb_2_1_FRAMING_ERR), .B(\data_out[4] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[4] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[5]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[5] ), 
        .D(\rx_byte[5] ), .Y(\NxtPrdata_5_am_0[5] ));
    SLE \controlReg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[5]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[0]  (.A(
        CoreUARTapb_2_1_TXRDY), .B(\data_out[0] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[0] ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[2]  (.A(
        \controlReg2[2]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[2]_net_1 ), .Y(\NxtPrdata_5_bm[2]_net_1 ));
    SLE \controlReg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[7]_net_1 ));
    SLE \iPRDATA[1]  (.D(\NxtPrdata[1] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[1]));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[6]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[6] ), 
        .D(\rx_byte[6] ), .Y(\NxtPrdata_5_am_1[6] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[7]  (.A(
        \controlReg2[7]_net_1 ), .B(\controlReg1[7]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[7] ));
    SLE \controlReg2[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[4]_net_1 ));
    SLE \iPRDATA[4]  (.D(\NxtPrdata[4] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[4]));
    VCC VCC (.Y(VCC_net_1));
    SLE \iPRDATA[3]  (.D(\NxtPrdata[3] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[3]));
    SLE \controlReg2[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[6]_net_1 ));
    SLE \controlReg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[3]_net_1 ));
    CFG4 #( .INIT(16'hC0A0) )  \NxtPrdata_5_0_a2[3]  (.A(
        \controlReg1[3]_net_1 ), .B(\controlReg2[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_606));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[4]  (.A(
        \controlReg2[4]_net_1 ), .B(\controlReg1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[4] ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[5]  (.A(
        \controlReg2[5]_net_1 ), .B(\controlReg1[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_0[5] ));
    SLE \controlReg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[0]  (.A(
        \controlReg2[0]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[0]_net_1 ), .Y(\NxtPrdata_5_bm_0[0] ));
    SLE \controlReg2[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[3]_net_1 ));
    SLE \controlReg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[2]_net_1 ));
    SLE \controlReg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[4]_net_1 ));
    SLE \iPRDATA[5]  (.D(\NxtPrdata[5] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[5]));
    SLE \iPRDATA[7]  (.D(\NxtPrdata[7] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[7]));
    CFG4 #( .INIT(16'hFFEC) )  \NxtPrdata_5_0[3]  (.A(\data_out[3] ), 
        .B(N_606), .C(N_367), .D(N_608), .Y(\NxtPrdata[3] ));
    SLE \controlReg2[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24_0_a2  (.A(
        CoreAPB3_0_APBmslave3_PSELx), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(controlReg24));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[6]  (.A(
        \controlReg2[6]_net_1 ), .B(\controlReg1[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm_1[6] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[4] ), .C(
        \NxtPrdata_5_am_0[4] ), .Y(\NxtPrdata[4] ));
    SLE \controlReg2[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[7]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[1]_net_1 ), 
        .C(\NxtPrdata_5_am[1]_net_1 ), .Y(\NxtPrdata[1] ));
    SLE \iPRDATA[2]  (.D(\NxtPrdata[2] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[2]));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[0] ), .C(
        \NxtPrdata_5_am_0[0] ), .Y(\NxtPrdata[0] ));
    SLE \controlReg2[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[5]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[1]  (.A(
        CoreUARTapb_2_1_RXRDY), .B(\data_out[1] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[1]_net_1 ));
    SLE \controlReg2[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[2]_net_1 ));
    SLE \iPRDATA[6]  (.D(\NxtPrdata[6] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[6]));
    SLE \iPRDATA[0]  (.D(\NxtPrdata[0] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave3_PRDATA[0]));
    mss_sb_CoreUARTapb_2_1_COREUART_1s_1s_0s_15s_0s uUART (
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .data_out({\data_out[4] , 
        \data_out[3] , \data_out[2] , \data_out[1] , \data_out[0] }), 
        .controlReg1({\controlReg1[7]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[5]_net_1 , \controlReg1[4]_net_1 , 
        \controlReg1[3]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[0]_net_1 }), .controlReg2({
        \controlReg2[7]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[1]_net_1 , \controlReg2[0]_net_1 }), 
        .rx_dout_reg_5(\rx_dout_reg[5] ), .rx_dout_reg_6(
        \rx_dout_reg[6] ), .rx_dout_reg_7(\rx_dout_reg[7] ), 
        .rx_byte_7(\rx_byte[7] ), .rx_byte_6(\rx_byte[6] ), .rx_byte_5(
        \rx_byte[5] ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreUARTapb_2_1_OVERFLOW(CoreUARTapb_2_1_OVERFLOW), 
        .CoreUARTapb_2_1_RXRDY(CoreUARTapb_2_1_RXRDY), .N_669(N_669), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreUARTapb_2_1_PARITY_ERR(CoreUARTapb_2_1_PARITY_ERR), 
        .N_367(N_367), .clear_overflow_0_a2_0_0(
        clear_overflow_0_a2_0_0), .GPS_RX_c(GPS_RX_c), 
        .CoreUARTapb_2_1_TXRDY(CoreUARTapb_2_1_TXRDY), .GPS_TX_c(
        GPS_TX_c), .CoreUARTapb_2_1_FRAMING_ERR(
        CoreUARTapb_2_1_FRAMING_ERR));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[7] ), .C(
        \NxtPrdata_5_am_0[7] ), .Y(\NxtPrdata[7] ));
    CFG2 #( .INIT(4'h4) )  \NxtPrdata_5_0_a2_2[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_425));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[2]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(\data_out[2] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[2]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \NxtPrdata_5_0_a2_1[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(N_425), .C(
        CoreUARTapb_2_1_OVERFLOW), .Y(N_608));
    SLE \controlReg2[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[0]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[2]_net_1 ), 
        .C(\NxtPrdata_5_am[2]_net_1 ), .Y(\NxtPrdata[2] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_1[6] ), .C(
        \NxtPrdata_5_am_1[6] ), .Y(\NxtPrdata[6] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[7]  (.A(
        CoreUARTapb_2_1_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[7] ), 
        .D(\rx_byte[7] ), .Y(\NxtPrdata_5_am_0[7] ));
    SLE \controlReg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[1]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \p_CtrlReg1Seq.controlReg14_0_a2  (.A(
        CoreAPB3_0_APBmslave3_PSELx), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(controlReg14));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[1]  (.A(
        \controlReg2[1]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[1]_net_1 ), .Y(\NxtPrdata_5_bm[1]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  un1_NxtPrdata23_i_a2 (.A(
        CoreAPB3_0_APBmslave0_PWRITE), .B(
        CoreAPB3_0_APBmslave0_PENABLE), .C(
        psh_negedge_reg_1_sqmuxa_6_2), .D(CoreAPB3_0_APBmslave3_PSELx), 
        .Y(un1_NxtPrdata23_i_a2_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[5] ), .C(
        \NxtPrdata_5_am_0[5] ), .Y(\NxtPrdata[5] ));
    SLE \controlReg1[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[0]_net_1 ));
    
endmodule


module pwm_gen_8s_16s_0(
       PWM_c,
       period_cnt,
       pwm_negedge_reg,
       pwm_enable_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST
    );
output [8:1] PWM_c;
input  [15:0] period_cnt;
input  [128:1] pwm_negedge_reg;
input  [8:1] pwm_enable_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;

    wire VCC_net_1, \PWM_int_108[8] , \un1_pwm_enable_reg_i_0[0] , 
        GND_net_1, N_509_i_0, \un1_pwm_enable_reg_1_i_0[0]_net_1 , 
        \PWM_int_80[6] , \un1_pwm_enable_reg_2_i_0[0] , N_26_i_0, N_62, 
        \PWM_int_52[4] , \un1_pwm_enable_reg_4_i_0[0] , N_508_i_0, 
        \un1_pwm_enable_reg_5_i_0[0]_net_1 , N_31_i_0, N_13, N_28_i_0, 
        \un1_pwm_enable_reg_7_0_a4_i[0]_net_1 , 
        \un1_period_cnt_1_0_data_tmp[0] , 
        \un1_period_cnt_1_0_data_tmp[1] , 
        \un1_period_cnt_1_0_data_tmp[2] , 
        \un1_period_cnt_1_0_data_tmp[3] , 
        \un1_period_cnt_1_0_data_tmp[4] , 
        \un1_period_cnt_1_0_data_tmp[5] , 
        \un1_period_cnt_1_0_data_tmp[6] , un1_period_cnt_1, 
        \un1_period_cnt_1_0_data_tmp_0[0] , 
        \un1_period_cnt_1_0_data_tmp_0[1] , 
        \un1_period_cnt_1_0_data_tmp_0[2] , 
        \un1_period_cnt_1_0_data_tmp_0[3] , 
        \un1_period_cnt_1_0_data_tmp_0[4] , 
        \un1_period_cnt_1_0_data_tmp_0[5] , 
        \un1_period_cnt_1_0_data_tmp_0[6] , un1_period_cnt_1_0, 
        \un1_period_cnt_1_0_data_tmp_1[0] , 
        \un1_period_cnt_1_0_data_tmp_1[1] , 
        \un1_period_cnt_1_0_data_tmp_1[2] , 
        \un1_period_cnt_1_0_data_tmp_1[3] , 
        \un1_period_cnt_1_0_data_tmp_1[4] , 
        \un1_period_cnt_1_0_data_tmp_1[5] , 
        \un1_period_cnt_1_0_data_tmp_1[6] , un1_period_cnt_1_1, 
        \un1_period_cnt_1_0_data_tmp_2[0] , 
        \un1_period_cnt_1_0_data_tmp_2[1] , 
        \un1_period_cnt_1_0_data_tmp_2[2] , 
        \un1_period_cnt_1_0_data_tmp_2[3] , 
        \un1_period_cnt_1_0_data_tmp_2[4] , 
        \un1_period_cnt_1_0_data_tmp_2[5] , 
        \un1_period_cnt_1_0_data_tmp_2[6] , un1_period_cnt_1_2, 
        \un1_period_cnt_1_0_data_tmp_3[0] , 
        \un1_period_cnt_1_0_data_tmp_3[1] , 
        \un1_period_cnt_1_0_data_tmp_3[2] , 
        \un1_period_cnt_1_0_data_tmp_3[3] , 
        \un1_period_cnt_1_0_data_tmp_3[4] , 
        \un1_period_cnt_1_0_data_tmp_3[5] , 
        \un1_period_cnt_1_0_data_tmp_3[6] , un1_period_cnt_1_3, 
        \un1_period_cnt_1_0_data_tmp_4[0] , 
        \un1_period_cnt_1_0_data_tmp_4[1] , 
        \un1_period_cnt_1_0_data_tmp_4[2] , 
        \un1_period_cnt_1_0_data_tmp_4[3] , 
        \un1_period_cnt_1_0_data_tmp_4[4] , 
        \un1_period_cnt_1_0_data_tmp_4[5] , 
        \un1_period_cnt_1_0_data_tmp_4[6] , un1_period_cnt_1_4, 
        \un1_period_cnt_1_0_data_tmp_5[0] , 
        \un1_period_cnt_1_0_data_tmp_5[1] , 
        \un1_period_cnt_1_0_data_tmp_5[2] , 
        \un1_period_cnt_1_0_data_tmp_5[3] , 
        \un1_period_cnt_1_0_data_tmp_5[4] , 
        \un1_period_cnt_1_0_data_tmp_5[5] , 
        \un1_period_cnt_1_0_data_tmp_5[6] , un1_period_cnt_1_5, 
        \un1_period_cnt_1_1_data_tmp[0] , 
        \un1_period_cnt_1_1_data_tmp[1] , 
        \un1_period_cnt_1_1_data_tmp[2] , 
        \un1_period_cnt_1_1_data_tmp[3] , 
        \un1_period_cnt_1_1_data_tmp[4] , 
        \un1_period_cnt_1_1_data_tmp[5] , 
        \un1_period_cnt_1_1_data_tmp[6] , un1_period_cnt_1_6, 
        \PWM_int_108_f1_2[8] , \PWM_int_94_f0_i_a2_2[7] , 
        \PWM_int_10_f0_i_0_a2_2[1] , \PWM_int_52_f1_2[4] , 
        \PWM_int_80_f1_2[6] , \PWM_int_38_f0_i_a2_2[3] , 
        \PWM_int_66_f0_i_0_a2_2[5] , \PWM_int_24_f0_i_0_a2_2[2] , 
        \PWM_int_108_f1_11[8] , \PWM_int_108_f1_10[8] , 
        \PWM_int_108_f1_8[8] , \PWM_int_24_f0_i_0_o2_11[2] , 
        \PWM_int_24_f0_i_0_o2_10[2] , \PWM_int_24_f0_i_0_o2_9[2] , 
        \PWM_int_24_f0_i_0_o2_8[2] , \PWM_int_94_f0_i_a2_11[7] , 
        \PWM_int_94_f0_i_a2_10[7] , \PWM_int_94_f0_i_a2_8[7] , 
        \PWM_int_10_f0_i_0_a2_11[1] , \PWM_int_10_f0_i_0_a2_10[1] , 
        \PWM_int_10_f0_i_0_a2_8[1] , \PWM_int_52_f1_11[4] , 
        \PWM_int_52_f1_10[4] , \PWM_int_52_f1_8[4] , 
        \PWM_int_80_f1_11[6] , \PWM_int_80_f1_10[6] , 
        \PWM_int_80_f1_8[6] , \PWM_int_38_f0_i_a2_11[3] , 
        \PWM_int_38_f0_i_a2_10[3] , \PWM_int_38_f0_i_a2_8[3] , 
        \PWM_int_66_f0_i_0_a2_11[5] , \PWM_int_66_f0_i_0_a2_10[5] , 
        \PWM_int_66_f0_i_0_a2_8[5] , \PWM_int_24_f0_i_0_a2_11[2] , 
        \PWM_int_24_f0_i_0_a2_10[2] , \PWM_int_24_f0_i_0_a2_8[2] , 
        \PWM_int_108_f1_13[8] , \PWM_int_94_f0_i_a2_13[7] , 
        \PWM_int_10_f0_i_0_a2_13[1] , \PWM_int_52_f1_13[4] , 
        \PWM_int_80_f1_13[6] , \PWM_int_38_f0_i_a2_13[3] , 
        \PWM_int_66_f0_i_0_a2_13[5] , \PWM_int_24_f0_i_0_a2_13[2] , 
        \PWM_int_108_f1_14[8] , \PWM_int_94_f0_i_a2_14[7] , 
        \PWM_int_10_f0_i_0_a2_14[1] , \PWM_int_52_f1_14[4] , 
        \PWM_int_80_f1_14[6] , \PWM_int_38_f0_i_a2_14[3] , 
        \PWM_int_66_f0_i_0_a2_14[5] , \PWM_int_24_f0_i_0_a2_14[2] , 
        N_218;
    
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[42]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[41]), .FCI(\un1_period_cnt_1_0_data_tmp_4[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_4[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_14[6]  (.A(
        pwm_negedge_reg[92]), .B(pwm_negedge_reg[91]), .C(
        \PWM_int_80_f1_11[6] ), .D(\PWM_int_80_f1_8[6] ), .Y(
        \PWM_int_80_f1_14[6] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_11[2]  
        (.A(pwm_negedge_reg[29]), .B(pwm_negedge_reg[21]), .C(
        pwm_negedge_reg[18]), .D(pwm_negedge_reg[17]), .Y(
        \PWM_int_24_f0_i_0_a2_11[2] ));
    SLE \PWM_output_generation[1].genblk1.PWM_int[1]  (.D(N_28_i_0), 
        .CLK(GL0_INST), .EN(\un1_pwm_enable_reg_7_0_a4_i[0]_net_1 ), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[1]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[120]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[119]), .FCI(
        \un1_period_cnt_1_0_data_tmp[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_10[4]  (.A(
        pwm_negedge_reg[60]), .B(pwm_negedge_reg[59]), .C(
        pwm_negedge_reg[58]), .D(pwm_negedge_reg[57]), .Y(
        \PWM_int_52_f1_10[4] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_14[8]  (.A(
        pwm_negedge_reg[115]), .B(pwm_negedge_reg[114]), .C(
        \PWM_int_108_f1_11[8] ), .D(\PWM_int_108_f1_8[8] ), .Y(
        \PWM_int_108_f1_14[8] ));
    CFG4 #( .INIT(16'h00A8) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f0[4]  (.A(
        pwm_enable_reg[4]), .B(\PWM_int_52_f1_13[4] ), .C(
        \PWM_int_52_f1_14[4] ), .D(N_218), .Y(\PWM_int_52[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[40]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[39]), .FCI(\un1_period_cnt_1_0_data_tmp_4[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_4[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_o2_10[2]  
        (.A(period_cnt[10]), .B(period_cnt[6]), .C(period_cnt[5]), .D(
        period_cnt[4]), .Y(\PWM_int_24_f0_i_0_o2_10[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[102]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[101]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[98]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[97]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[0] ));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_2[6]  (.A(
        pwm_negedge_reg[85]), .B(pwm_negedge_reg[86]), .Y(
        \PWM_int_80_f1_2[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_1  (.A(
        pwm_negedge_reg[2]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[1]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_1_data_tmp[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[108]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[107]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[5] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_13[5]  
        (.A(pwm_negedge_reg[65]), .B(pwm_negedge_reg[66]), .C(
        \PWM_int_66_f0_i_0_a2_10[5] ), .D(\PWM_int_66_f0_i_0_a2_2[5] ), 
        .Y(\PWM_int_66_f0_i_0_a2_13[5] ));
    CFG3 #( .INIT(8'hDF) )  
        \PWM_output_generation[8].genblk1.PWM_int_RNO[8]  (.A(
        pwm_enable_reg[8]), .B(un1_period_cnt_1), .C(N_218), .Y(
        \un1_pwm_enable_reg_i_0[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_45  (.A(
        pwm_negedge_reg[16]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[15]), .FCI(\un1_period_cnt_1_1_data_tmp[6] )
        , .S(), .Y(), .FCO(un1_period_cnt_1_6));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_11[6]  (.A(
        pwm_negedge_reg[96]), .B(pwm_negedge_reg[95]), .C(
        pwm_negedge_reg[94]), .D(pwm_negedge_reg[93]), .Y(
        \PWM_int_80_f1_11[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_39  (.A(
        pwm_negedge_reg[4]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[3]), .FCI(\un1_period_cnt_1_1_data_tmp[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_15  (.A(
        pwm_negedge_reg[12]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[11]), .FCI(\un1_period_cnt_1_1_data_tmp[4] )
        , .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[62]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[61]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[6] ));
    SLE \PWM_output_generation[3].genblk1.PWM_int[3]  (.D(N_508_i_0), 
        .CLK(GL0_INST), .EN(\un1_pwm_enable_reg_5_i_0[0]_net_1 ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[3]));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_2[4]  (.A(
        pwm_negedge_reg[63]), .B(pwm_negedge_reg[64]), .Y(
        \PWM_int_52_f1_2[4] ));
    CFG4 #( .INIT(16'h002A) )  
        \PWM_output_generation[3].genblk1.PWM_int_RNO[3]  (.A(
        pwm_enable_reg[3]), .B(\PWM_int_38_f0_i_a2_13[3] ), .C(
        \PWM_int_38_f0_i_a2_14[3] ), .D(N_218), .Y(N_508_i_0));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_8[7]  (.A(
        pwm_negedge_reg[110]), .B(pwm_negedge_reg[102]), .C(PWM_c[7]), 
        .Y(\PWM_int_94_f0_i_a2_8[7] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_13[4]  (.A(
        pwm_negedge_reg[61]), .B(pwm_negedge_reg[62]), .C(
        \PWM_int_52_f1_10[4] ), .D(\PWM_int_52_f1_2[4] ), .Y(
        \PWM_int_52_f1_13[4] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_8[8]  (.A(
        pwm_negedge_reg[128]), .B(pwm_negedge_reg[113]), .C(PWM_c[8]), 
        .Y(\PWM_int_108_f1_8[8] ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_o2_9[2]  (
        .A(period_cnt[7]), .B(period_cnt[3]), .C(period_cnt[2]), .D(
        period_cnt[1]), .Y(\PWM_int_24_f0_i_0_o2_9[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[50]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[49]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[52]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[51]), .FCI(\un1_period_cnt_1_0_data_tmp_3[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[32]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[31]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_5));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_10[7]  (
        .A(pwm_negedge_reg[112]), .B(pwm_negedge_reg[111]), .C(
        pwm_negedge_reg[107]), .D(pwm_negedge_reg[98]), .Y(
        \PWM_int_94_f0_i_a2_10[7] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_13[8]  (.A(
        pwm_negedge_reg[126]), .B(pwm_negedge_reg[127]), .C(
        \PWM_int_108_f1_10[8] ), .D(\PWM_int_108_f1_2[8] ), .Y(
        \PWM_int_108_f1_13[8] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_10[3]  (
        .A(pwm_negedge_reg[36]), .B(pwm_negedge_reg[35]), .C(
        pwm_negedge_reg[34]), .D(pwm_negedge_reg[33]), .Y(
        \PWM_int_38_f0_i_a2_10[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[106]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[105]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[4] ));
    CFG2 #( .INIT(4'h1) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_2[2]  (
        .A(pwm_negedge_reg[20]), .B(pwm_negedge_reg[22]), .Y(
        \PWM_int_24_f0_i_0_a2_2[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[60]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[59]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_3[5] ));
    CFG4 #( .INIT(16'h002A) )  
        \PWM_output_generation[2].genblk1.PWM_int_RNO[2]  (.A(
        pwm_enable_reg[2]), .B(\PWM_int_24_f0_i_0_a2_13[2] ), .C(
        \PWM_int_24_f0_i_0_a2_14[2] ), .D(N_218), .Y(N_31_i_0));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[116]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[115]), .FCI(
        \un1_period_cnt_1_0_data_tmp[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[1] ));
    CFG3 #( .INIT(8'hDF) )  \un1_pwm_enable_reg_1_i_0[0]  (.A(
        pwm_enable_reg[7]), .B(un1_period_cnt_1_0), .C(N_218), .Y(
        \un1_pwm_enable_reg_1_i_0[0]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  \un1_pwm_enable_reg_5_i_0[0]  (.A(
        pwm_enable_reg[3]), .B(un1_period_cnt_1_4), .C(N_218), .Y(
        \un1_pwm_enable_reg_5_i_0[0]_net_1 ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[104]), .B(period_cnt[6]), .C(period_cnt[7]), 
        .D(pwm_negedge_reg[103]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[2] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[3] ));
    SLE \PWM_output_generation[2].genblk1.PWM_int[2]  (.D(N_31_i_0), 
        .CLK(GL0_INST), .EN(N_13), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[2]));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_11[7]  (
        .A(pwm_negedge_reg[109]), .B(pwm_negedge_reg[106]), .C(
        pwm_negedge_reg[105]), .D(pwm_negedge_reg[97]), .Y(
        \PWM_int_94_f0_i_a2_11[7] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[46]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[45]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[84]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[83]), .FCI(\un1_period_cnt_1_0_data_tmp_1[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_11[8]  (.A(
        pwm_negedge_reg[119]), .B(pwm_negedge_reg[118]), .C(
        pwm_negedge_reg[117]), .D(pwm_negedge_reg[116]), .Y(
        \PWM_int_108_f1_11[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_27  (.A(
        pwm_negedge_reg[10]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[9]), .FCI(\un1_period_cnt_1_1_data_tmp[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[4] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_11[5]  
        (.A(pwm_negedge_reg[80]), .B(pwm_negedge_reg[79]), .C(
        pwm_negedge_reg[70]), .D(pwm_negedge_reg[69]), .Y(
        \PWM_int_66_f0_i_0_a2_11[5] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_o2_11[2]  
        (.A(period_cnt[13]), .B(period_cnt[11]), .C(period_cnt[9]), .D(
        period_cnt[8]), .Y(\PWM_int_24_f0_i_0_o2_11[2] ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_o2_8[2]  (
        .A(period_cnt[15]), .B(period_cnt[14]), .C(period_cnt[12]), .D(
        period_cnt[0]), .Y(\PWM_int_24_f0_i_0_o2_8[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_11[4]  (.A(
        pwm_negedge_reg[52]), .B(pwm_negedge_reg[51]), .C(
        pwm_negedge_reg[50]), .D(pwm_negedge_reg[49]), .Y(
        \PWM_int_52_f1_11[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_33  (.A(
        pwm_negedge_reg[6]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[5]), .FCI(\un1_period_cnt_1_1_data_tmp[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[90]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[89]), .FCI(\un1_period_cnt_1_0_data_tmp_1[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[4] ));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_8[3]  (.A(
        pwm_negedge_reg[41]), .B(pwm_negedge_reg[40]), .C(PWM_c[3]), 
        .Y(\PWM_int_38_f0_i_a2_8[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_21  (.A(
        pwm_negedge_reg[8]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[7]), .FCI(\un1_period_cnt_1_1_data_tmp[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[36]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[35]), .FCI(\un1_period_cnt_1_0_data_tmp_4[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_4[1] ));
    SLE \PWM_output_generation[7].genblk1.PWM_int[7]  (.D(N_509_i_0), 
        .CLK(GL0_INST), .EN(\un1_pwm_enable_reg_1_i_0[0]_net_1 ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[7]));
    SLE \PWM_output_generation[6].genblk1.PWM_int[6]  (.D(
        \PWM_int_80[6] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_2_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[6]));
    CFG2 #( .INIT(4'hE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_2[8]  (.A(
        pwm_negedge_reg[124]), .B(pwm_negedge_reg[125]), .Y(
        \PWM_int_108_f1_2[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[88]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[87]), .FCI(\un1_period_cnt_1_0_data_tmp_1[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[3] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_11[1]  
        (.A(pwm_negedge_reg[13]), .B(pwm_negedge_reg[10]), .C(
        pwm_negedge_reg[9]), .D(pwm_negedge_reg[1]), .Y(
        \PWM_int_10_f0_i_0_a2_11[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[112]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[111]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_0));
    CFG4 #( .INIT(16'h00A8) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f0[6]  (.A(
        pwm_enable_reg[6]), .B(\PWM_int_80_f1_13[6] ), .C(
        \PWM_int_80_f1_14[6] ), .D(N_218), .Y(\PWM_int_80[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[54]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[53]), .FCI(\un1_period_cnt_1_0_data_tmp_3[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[34]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[33]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[0] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_13[1]  
        (.A(pwm_negedge_reg[14]), .B(pwm_negedge_reg[16]), .C(
        \PWM_int_10_f0_i_0_a2_10[1] ), .D(\PWM_int_10_f0_i_0_a2_2[1] ), 
        .Y(\PWM_int_10_f0_i_0_a2_13[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[1].genblk1.un1_period_cnt_1_1_I_9  (.A(
        pwm_negedge_reg[14]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[13]), .FCI(\un1_period_cnt_1_1_data_tmp[5] )
        , .S(), .Y(), .FCO(\un1_period_cnt_1_1_data_tmp[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[18]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[17]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_13[6]  (.A(
        pwm_negedge_reg[87]), .B(pwm_negedge_reg[88]), .C(
        \PWM_int_80_f1_10[6] ), .D(\PWM_int_80_f1_2[6] ), .Y(
        \PWM_int_80_f1_13[6] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_8[4]  (.A(
        pwm_negedge_reg[54]), .B(pwm_negedge_reg[53]), .C(PWM_c[4]), 
        .Y(\PWM_int_52_f1_8[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[118]), .B(period_cnt[4]), .C(period_cnt[5]), 
        .D(pwm_negedge_reg[117]), .FCI(
        \un1_period_cnt_1_0_data_tmp[1] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[44]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[43]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_4[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[20]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[19]), .FCI(\un1_period_cnt_1_0_data_tmp_5[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_5[1] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_10[2]  
        (.A(pwm_negedge_reg[32]), .B(pwm_negedge_reg[31]), .C(
        pwm_negedge_reg[27]), .D(pwm_negedge_reg[25]), .Y(
        \PWM_int_24_f0_i_0_a2_10[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[28]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[27]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[5] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_14[7]  (
        .A(pwm_negedge_reg[108]), .B(pwm_negedge_reg[101]), .C(
        \PWM_int_94_f0_i_a2_11[7] ), .D(\PWM_int_94_f0_i_a2_8[7] ), .Y(
        \PWM_int_94_f0_i_a2_14[7] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[86]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[85]), .FCI(\un1_period_cnt_1_0_data_tmp_1[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_1[2] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_14[3]  (
        .A(pwm_negedge_reg[45]), .B(pwm_negedge_reg[39]), .C(
        \PWM_int_38_f0_i_a2_11[3] ), .D(\PWM_int_38_f0_i_a2_8[3] ), .Y(
        \PWM_int_38_f0_i_a2_14[3] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[66]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[65]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[110]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[109]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[6] ));
    CFG4 #( .INIT(16'h002A) )  
        \PWM_output_generation[1].genblk1.PWM_int_RNO[1]  (.A(
        pwm_enable_reg[1]), .B(\PWM_int_10_f0_i_0_a2_13[1] ), .C(
        \PWM_int_10_f0_i_0_a2_14[1] ), .D(N_218), .Y(N_28_i_0));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[96]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[95]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_1));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_14[1]  
        (.A(pwm_negedge_reg[12]), .B(pwm_negedge_reg[11]), .C(
        \PWM_int_10_f0_i_0_a2_11[1] ), .D(\PWM_int_10_f0_i_0_a2_8[1] ), 
        .Y(\PWM_int_10_f0_i_0_a2_14[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[68]), .B(period_cnt[2]), .C(period_cnt[3]), .D(
        pwm_negedge_reg[67]), .FCI(\un1_period_cnt_1_0_data_tmp_2[0] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[1] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_11[3]  (
        .A(pwm_negedge_reg[48]), .B(pwm_negedge_reg[47]), .C(
        pwm_negedge_reg[38]), .D(pwm_negedge_reg[37]), .Y(
        \PWM_int_38_f0_i_a2_11[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_o2[2]  (.A(
        \PWM_int_24_f0_i_0_o2_11[2] ), .B(\PWM_int_24_f0_i_0_o2_10[2] )
        , .C(\PWM_int_24_f0_i_0_o2_9[2] ), .D(
        \PWM_int_24_f0_i_0_o2_8[2] ), .Y(N_218));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[76]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[75]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[5] ));
    CFG3 #( .INIT(8'hEF) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_8[6]  (.A(
        pwm_negedge_reg[90]), .B(pwm_negedge_reg[89]), .C(PWM_c[6]), 
        .Y(\PWM_int_80_f1_8[6] ));
    SLE \PWM_output_generation[5].genblk1.PWM_int[5]  (.D(N_26_i_0), 
        .CLK(GL0_INST), .EN(N_62), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[5]));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[38]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[37]), .FCI(\un1_period_cnt_1_0_data_tmp_4[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_4[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[4].genblk1.PWM_int_52_f1_14[4]  (.A(
        pwm_negedge_reg[56]), .B(pwm_negedge_reg[55]), .C(
        \PWM_int_52_f1_11[4] ), .D(\PWM_int_52_f1_8[4] ), .Y(
        \PWM_int_52_f1_14[4] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_13[3]  (
        .A(pwm_negedge_reg[42]), .B(pwm_negedge_reg[44]), .C(
        \PWM_int_38_f0_i_a2_10[3] ), .D(\PWM_int_38_f0_i_a2_2[3] ), .Y(
        \PWM_int_38_f0_i_a2_13[3] ));
    CFG4 #( .INIT(16'h002A) )  
        \PWM_output_generation[5].genblk1.PWM_int_RNO[5]  (.A(
        pwm_enable_reg[5]), .B(\PWM_int_66_f0_i_0_a2_13[5] ), .C(
        \PWM_int_66_f0_i_0_a2_14[5] ), .D(N_218), .Y(N_26_i_0));
    CFG3 #( .INIT(8'hDF) )  \un1_pwm_enable_reg_6_i_0_0[0]  (.A(
        pwm_enable_reg[2]), .B(un1_period_cnt_1_5), .C(N_218), .Y(N_13)
        );
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[114]), .B(period_cnt[0]), .C(period_cnt[1]), 
        .D(pwm_negedge_reg[113]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[0] ));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_8[1]  (
        .A(pwm_negedge_reg[7]), .B(pwm_negedge_reg[6]), .C(PWM_c[1]), 
        .Y(\PWM_int_10_f0_i_0_a2_8[1] ));
    CFG2 #( .INIT(4'h1) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_2[1]  (
        .A(pwm_negedge_reg[3]), .B(pwm_negedge_reg[8]), .Y(
        \PWM_int_10_f0_i_0_a2_2[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[124]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[123]), .FCI(
        \un1_period_cnt_1_0_data_tmp[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[3].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[48]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[47]), .FCI(
        \un1_period_cnt_1_0_data_tmp_4[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_4));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[30]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[29]), .FCI(
        \un1_period_cnt_1_0_data_tmp_5[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_5[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[128]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[127]), .FCI(
        \un1_period_cnt_1_0_data_tmp[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[6].genblk1.PWM_int_80_f1_10[6]  (.A(
        pwm_negedge_reg[84]), .B(pwm_negedge_reg[83]), .C(
        pwm_negedge_reg[82]), .D(pwm_negedge_reg[81]), .Y(
        \PWM_int_80_f1_10[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_1  (.A(
        pwm_negedge_reg[82]), .B(period_cnt[0]), .C(period_cnt[1]), .D(
        pwm_negedge_reg[81]), .FCI(VCC_net_1), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[0] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[22]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[21]), .FCI(\un1_period_cnt_1_0_data_tmp_5[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_5[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[74]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[73]), .FCI(\un1_period_cnt_1_0_data_tmp_2[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_15  (.A(
        pwm_negedge_reg[92]), .B(period_cnt[10]), .C(period_cnt[11]), 
        .D(pwm_negedge_reg[91]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[4] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[5] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[7].genblk1.un1_period_cnt_1_0_I_39  (.A(
        pwm_negedge_reg[100]), .B(period_cnt[2]), .C(period_cnt[3]), 
        .D(pwm_negedge_reg[99]), .FCI(
        \un1_period_cnt_1_0_data_tmp_0[0] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_0[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[58]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[57]), .FCI(\un1_period_cnt_1_0_data_tmp_3[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[4] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[78]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[77]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_2[6] ));
    CFG2 #( .INIT(4'h1) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_2[5]  (
        .A(pwm_negedge_reg[67]), .B(pwm_negedge_reg[68]), .Y(
        \PWM_int_66_f0_i_0_a2_2[5] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_14[5]  
        (.A(pwm_negedge_reg[77]), .B(pwm_negedge_reg[71]), .C(
        \PWM_int_66_f0_i_0_a2_11[5] ), .D(\PWM_int_66_f0_i_0_a2_8[5] ), 
        .Y(\PWM_int_66_f0_i_0_a2_14[5] ));
    CFG4 #( .INIT(16'h00A8) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f0[8]  (.A(
        pwm_enable_reg[8]), .B(\PWM_int_108_f1_13[8] ), .C(
        \PWM_int_108_f1_14[8] ), .D(N_218), .Y(\PWM_int_108[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[72]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[71]), .FCI(\un1_period_cnt_1_0_data_tmp_2[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \PWM_output_generation[8].genblk1.PWM_int_108_f1_10[8]  (.A(
        pwm_negedge_reg[123]), .B(pwm_negedge_reg[122]), .C(
        pwm_negedge_reg[121]), .D(pwm_negedge_reg[120]), .Y(
        \PWM_int_108_f1_10[8] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_33  (.A(
        pwm_negedge_reg[70]), .B(period_cnt[4]), .C(period_cnt[5]), .D(
        pwm_negedge_reg[69]), .FCI(\un1_period_cnt_1_0_data_tmp_2[1] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_2[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[126]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[125]), .FCI(
        \un1_period_cnt_1_0_data_tmp[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[6] ));
    CFG3 #( .INIT(8'hDF) )  \un1_pwm_enable_reg_7_0_a4_i[0]  (.A(
        pwm_enable_reg[1]), .B(un1_period_cnt_1_6), .C(N_218), .Y(
        \un1_pwm_enable_reg_7_0_a4_i[0]_net_1 ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[26]), .B(period_cnt[8]), .C(period_cnt[9]), .D(
        pwm_negedge_reg[25]), .FCI(\un1_period_cnt_1_0_data_tmp_5[3] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_5[4] ));
    SLE \PWM_output_generation[4].genblk1.PWM_int[4]  (.D(
        \PWM_int_52[4] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_4_i_0[0] ), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(PWM_c[4]));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_10[5]  
        (.A(pwm_negedge_reg[78]), .B(pwm_negedge_reg[75]), .C(
        pwm_negedge_reg[74]), .D(pwm_negedge_reg[73]), .Y(
        \PWM_int_66_f0_i_0_a2_10[5] ));
    CFG3 #( .INIT(8'hDF) )  
        \PWM_output_generation[4].genblk1.PWM_int_RNO[4]  (.A(
        pwm_enable_reg[4]), .B(un1_period_cnt_1_3), .C(N_218), .Y(
        \un1_pwm_enable_reg_4_i_0[0] ));
    CFG2 #( .INIT(4'h1) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_2[7]  (.A(
        pwm_negedge_reg[99]), .B(pwm_negedge_reg[100]), .Y(
        \PWM_int_94_f0_i_a2_2[7] ));
    CFG4 #( .INIT(16'h0001) )  
        \PWM_output_generation[1].genblk1.PWM_int_10_f0_i_0_a2_10[1]  
        (.A(pwm_negedge_reg[15]), .B(pwm_negedge_reg[5]), .C(
        pwm_negedge_reg[4]), .D(pwm_negedge_reg[2]), .Y(
        \PWM_int_10_f0_i_0_a2_10[1] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[5].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[80]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[79]), .FCI(
        \un1_period_cnt_1_0_data_tmp_2[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_2));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[56]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[55]), .FCI(\un1_period_cnt_1_0_data_tmp_3[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_3[3] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_13[2]  
        (.A(pwm_negedge_reg[19]), .B(pwm_negedge_reg[30]), .C(
        \PWM_int_24_f0_i_0_a2_10[2] ), .D(\PWM_int_24_f0_i_0_a2_2[2] ), 
        .Y(\PWM_int_24_f0_i_0_a2_13[2] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[7].genblk1.PWM_int_94_f0_i_a2_13[7]  (
        .A(pwm_negedge_reg[103]), .B(pwm_negedge_reg[104]), .C(
        \PWM_int_94_f0_i_a2_10[7] ), .D(\PWM_int_94_f0_i_a2_2[7] ), .Y(
        \PWM_int_94_f0_i_a2_13[7] ));
    CFG4 #( .INIT(16'h002A) )  
        \PWM_output_generation[7].genblk1.PWM_int_RNO[7]  (.A(
        pwm_enable_reg[7]), .B(\PWM_int_94_f0_i_a2_13[7] ), .C(
        \PWM_int_94_f0_i_a2_14[7] ), .D(N_218), .Y(N_509_i_0));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[6].genblk1.un1_period_cnt_1_0_I_9  (.A(
        pwm_negedge_reg[94]), .B(period_cnt[12]), .C(period_cnt[13]), 
        .D(pwm_negedge_reg[93]), .FCI(
        \un1_period_cnt_1_0_data_tmp_1[5] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp_1[6] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[4].genblk1.un1_period_cnt_1_0_I_45  (.A(
        pwm_negedge_reg[64]), .B(period_cnt[14]), .C(period_cnt[15]), 
        .D(pwm_negedge_reg[63]), .FCI(
        \un1_period_cnt_1_0_data_tmp_3[6] ), .S(), .Y(), .FCO(
        un1_period_cnt_1_3));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[2].genblk1.un1_period_cnt_1_0_I_21  (.A(
        pwm_negedge_reg[24]), .B(period_cnt[6]), .C(period_cnt[7]), .D(
        pwm_negedge_reg[23]), .FCI(\un1_period_cnt_1_0_data_tmp_5[2] ), 
        .S(), .Y(), .FCO(\un1_period_cnt_1_0_data_tmp_5[3] ));
    CFG4 #( .INIT(16'h1000) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_14[2]  
        (.A(pwm_negedge_reg[28]), .B(pwm_negedge_reg[26]), .C(
        \PWM_int_24_f0_i_0_a2_11[2] ), .D(\PWM_int_24_f0_i_0_a2_8[2] ), 
        .Y(\PWM_int_24_f0_i_0_a2_14[2] ));
    CFG3 #( .INIT(8'hDF) )  \un1_pwm_enable_reg_3_0_a4_i[0]  (.A(
        pwm_enable_reg[5]), .B(un1_period_cnt_1_2), .C(N_218), .Y(N_62)
        );
    SLE \PWM_output_generation[8].genblk1.PWM_int[8]  (.D(
        \PWM_int_108[8] ), .CLK(GL0_INST), .EN(
        \un1_pwm_enable_reg_i_0[0] ), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(PWM_c[8]));
    CFG2 #( .INIT(4'h1) )  
        \PWM_output_generation[3].genblk1.PWM_int_38_f0_i_a2_2[3]  (.A(
        pwm_negedge_reg[43]), .B(pwm_negedge_reg[46]), .Y(
        \PWM_int_38_f0_i_a2_2[3] ));
    CFG3 #( .INIT(8'hDF) )  
        \PWM_output_generation[6].genblk1.PWM_int_RNO[6]  (.A(
        pwm_enable_reg[6]), .B(un1_period_cnt_1_1), .C(N_218), .Y(
        \un1_pwm_enable_reg_2_i_0[0] ));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[2].genblk1.PWM_int_24_f0_i_0_a2_8[2]  (
        .A(pwm_negedge_reg[24]), .B(pwm_negedge_reg[23]), .C(PWM_c[2]), 
        .Y(\PWM_int_24_f0_i_0_a2_8[2] ));
    ARI1 #( .INIT(20'h48421) )  
        \PWM_output_generation[8].genblk1.un1_period_cnt_1_0_I_27  (.A(
        pwm_negedge_reg[122]), .B(period_cnt[8]), .C(period_cnt[9]), 
        .D(pwm_negedge_reg[121]), .FCI(
        \un1_period_cnt_1_0_data_tmp[3] ), .S(), .Y(), .FCO(
        \un1_period_cnt_1_0_data_tmp[4] ));
    CFG3 #( .INIT(8'h10) )  
        \PWM_output_generation[5].genblk1.PWM_int_66_f0_i_0_a2_8[5]  (
        .A(pwm_negedge_reg[76]), .B(pwm_negedge_reg[72]), .C(PWM_c[5]), 
        .Y(\PWM_int_66_f0_i_0_a2_8[5] ));
    
endmodule


module timebase_16s(
       period_cnt,
       period_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST
    );
output [15:0] period_cnt;
input  [15:0] period_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;

    wire VCC_net_1, \period_cnt_s[0] , GND_net_1, \period_cnt_s[1] , 
        \period_cnt_s[2] , \period_cnt_s[3] , \period_cnt_s[4] , 
        \period_cnt_s[5] , \period_cnt_s[6] , \period_cnt_s[7] , 
        \period_cnt_s[8] , \period_cnt_s[9] , \period_cnt_s[10] , 
        \period_cnt_s[11] , \period_cnt_s[12] , \period_cnt_s[13] , 
        \period_cnt_s[14] , \period_cnt_s[15]_net_1 , 
        un1_period_cnt_cry_0_net_1, un1_period_cnt_cry_1_net_1, 
        un1_period_cnt_cry_2_net_1, un1_period_cnt_cry_3_net_1, 
        un1_period_cnt_cry_4_net_1, un1_period_cnt_cry_5_net_1, 
        un1_period_cnt_cry_6_net_1, un1_period_cnt_cry_7_net_1, 
        un1_period_cnt_cry_8_net_1, un1_period_cnt_cry_9_net_1, 
        un1_period_cnt_cry_10_net_1, un1_period_cnt_cry_11_net_1, 
        un1_period_cnt_cry_12_net_1, un1_period_cnt_cry_13_net_1, 
        un1_period_cnt_cry_14_net_1, period_cnt_net_1, 
        period_cnt_s_316_FCO, \period_cnt_cry[0]_net_1 , 
        \period_cnt_cry[1]_net_1 , \period_cnt_cry[2]_net_1 , 
        \period_cnt_cry[3]_net_1 , \period_cnt_cry[4]_net_1 , 
        \period_cnt_cry[5]_net_1 , \period_cnt_cry[6]_net_1 , 
        \period_cnt_cry[7]_net_1 , \period_cnt_cry[8]_net_1 , 
        \period_cnt_cry[9]_net_1 , \period_cnt_cry[10]_net_1 , 
        \period_cnt_cry[11]_net_1 , \period_cnt_cry[12]_net_1 , 
        \period_cnt_cry[13]_net_1 , \period_cnt_cry[14]_net_1 ;
    
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_9 (.A(period_reg[9])
        , .B(period_cnt[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_8_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_9_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_2 (.A(period_reg[2])
        , .B(period_cnt[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_1_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_2_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[14]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[14]), .D(GND_net_1), .FCI(
        \period_cnt_cry[13]_net_1 ), .S(\period_cnt_s[14] ), .Y(), 
        .FCO(\period_cnt_cry[14]_net_1 ));
    SLE \period_cnt[9]  (.D(\period_cnt_s[9] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[9]));
    SLE \period_cnt[6]  (.D(\period_cnt_s[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[6]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[0]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[0]), .D(GND_net_1), .FCI(
        period_cnt_s_316_FCO), .S(\period_cnt_s[0] ), .Y(), .FCO(
        \period_cnt_cry[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[8]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[8]), .D(GND_net_1), .FCI(
        \period_cnt_cry[7]_net_1 ), .S(\period_cnt_s[8] ), .Y(), .FCO(
        \period_cnt_cry[8]_net_1 ));
    SLE \period_cnt[14]  (.D(\period_cnt_s[14] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[14]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[11]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[11]), .D(GND_net_1), .FCI(
        \period_cnt_cry[10]_net_1 ), .S(\period_cnt_s[11] ), .Y(), 
        .FCO(\period_cnt_cry[11]_net_1 ));
    SLE \period_cnt[10]  (.D(\period_cnt_s[10] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[10]));
    SLE \period_cnt[0]  (.D(\period_cnt_s[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[0]));
    SLE \period_cnt[11]  (.D(\period_cnt_s[11] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[11]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_3 (.A(period_reg[3])
        , .B(period_cnt[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_2_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_3_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE \period_cnt[13]  (.D(\period_cnt_s[13] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[13]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[7]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[7]), .D(GND_net_1), .FCI(
        \period_cnt_cry[6]_net_1 ), .S(\period_cnt_s[7] ), .Y(), .FCO(
        \period_cnt_cry[7]_net_1 ));
    SLE \period_cnt[1]  (.D(\period_cnt_s[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[1]));
    SLE \period_cnt[7]  (.D(\period_cnt_s[7] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[7]));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[1]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[1]), .D(GND_net_1), .FCI(
        \period_cnt_cry[0]_net_1 ), .S(\period_cnt_s[1] ), .Y(), .FCO(
        \period_cnt_cry[1]_net_1 ));
    SLE \period_cnt[15]  (.D(\period_cnt_s[15]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(period_cnt[15]));
    SLE \period_cnt[2]  (.D(\period_cnt_s[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[2]));
    SLE \period_cnt[3]  (.D(\period_cnt_s[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[3]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_5 (.A(period_reg[5])
        , .B(period_cnt[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_4_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_5_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[9]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[9]), .D(GND_net_1), .FCI(
        \period_cnt_cry[8]_net_1 ), .S(\period_cnt_s[9] ), .Y(), .FCO(
        \period_cnt_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[2]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[2]), .D(GND_net_1), .FCI(
        \period_cnt_cry[1]_net_1 ), .S(\period_cnt_s[2] ), .Y(), .FCO(
        \period_cnt_cry[2]_net_1 ));
    SLE \period_cnt[5]  (.D(\period_cnt_s[5] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[5]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_11 (.A(
        period_reg[11]), .B(period_cnt[11]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_10_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_11_net_1));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[10]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[10]), .D(GND_net_1), .FCI(
        \period_cnt_cry[9]_net_1 ), .S(\period_cnt_s[10] ), .Y(), .FCO(
        \period_cnt_cry[10]_net_1 ));
    SLE \period_cnt[4]  (.D(\period_cnt_s[4] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[4]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_8 (.A(period_reg[8])
        , .B(period_cnt[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_7_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_8_net_1));
    SLE \period_cnt[8]  (.D(\period_cnt_s[8] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[8]));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_10 (.A(
        period_reg[10]), .B(period_cnt[10]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_9_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_10_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[12]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[12]), .D(GND_net_1), .FCI(
        \period_cnt_cry[11]_net_1 ), .S(\period_cnt_s[12] ), .Y(), 
        .FCO(\period_cnt_cry[12]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_4 (.A(period_reg[4])
        , .B(period_cnt[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_3_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_4_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_14 (.A(
        period_reg[14]), .B(period_cnt[14]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_13_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_14_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_7 (.A(period_reg[7])
        , .B(period_cnt[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_6_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_7_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_15 (.A(
        period_reg[15]), .B(period_cnt[15]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_14_net_1), .S(), .Y(), 
        .FCO(period_cnt_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[3]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[3]), .D(GND_net_1), .FCI(
        \period_cnt_cry[2]_net_1 ), .S(\period_cnt_s[3] ), .Y(), .FCO(
        \period_cnt_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[5]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[5]), .D(GND_net_1), .FCI(
        \period_cnt_cry[4]_net_1 ), .S(\period_cnt_s[5] ), .Y(), .FCO(
        \period_cnt_cry[5]_net_1 ));
    SLE \period_cnt[12]  (.D(\period_cnt_s[12] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        period_cnt[12]));
    ARI1 #( .INIT(20'h4AA00) )  period_cnt_s_316 (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(period_cnt_s_316_FCO));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_0 (.A(period_reg[0])
        , .B(period_cnt[0]), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(un1_period_cnt_cry_0_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[4]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[4]), .D(GND_net_1), .FCI(
        \period_cnt_cry[3]_net_1 ), .S(\period_cnt_s[4] ), .Y(), .FCO(
        \period_cnt_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_6 (.A(period_reg[6])
        , .B(period_cnt[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_5_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_6_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_12 (.A(
        period_reg[12]), .B(period_cnt[12]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_11_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_12_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_1 (.A(period_reg[1])
        , .B(period_cnt[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_0_net_1), .S(), .Y(), .FCO(
        un1_period_cnt_cry_1_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_s[15]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[15]), .D(GND_net_1), .FCI(
        \period_cnt_cry[14]_net_1 ), .S(\period_cnt_s[15]_net_1 ), .Y()
        , .FCO());
    ARI1 #( .INIT(20'h5AA55) )  un1_period_cnt_cry_13 (.A(
        period_reg[13]), .B(period_cnt[13]), .C(GND_net_1), .D(
        GND_net_1), .FCI(un1_period_cnt_cry_12_net_1), .S(), .Y(), 
        .FCO(un1_period_cnt_cry_13_net_1));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[13]  (.A(VCC_net_1), 
        .B(period_cnt_net_1), .C(period_cnt[13]), .D(GND_net_1), .FCI(
        \period_cnt_cry[12]_net_1 ), .S(\period_cnt_s[13] ), .Y(), 
        .FCO(\period_cnt_cry[13]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \period_cnt_cry[6]  (.A(VCC_net_1), .B(
        period_cnt_net_1), .C(period_cnt[6]), .D(GND_net_1), .FCI(
        \period_cnt_cry[5]_net_1 ), .S(\period_cnt_s[6] ), .Y(), .FCO(
        \period_cnt_cry[6]_net_1 ));
    
endmodule


module reg_if_Z5_layer0(
       CoreAPB3_0_APBmslave0_PWDATA,
       pwm_enable_reg,
       pwm_negedge_reg,
       period_reg,
       period_cnt,
       PRDATA_regif_0_0,
       CoreAPB3_0_APBmslave0_PADDR,
       PRDATA_regif_12_0,
       PRDATA_regif_9_i_1,
       PRDATA_regif_9_i_0_4,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_428,
       N_629,
       N_678,
       N_689,
       N_686,
       N_679,
       N_687,
       N_688,
       N_690,
       N_680,
       N_685,
       N_681,
       N_684,
       N_691,
       psh_enable_reg1_1_sqmuxa_0,
       N_528,
       psh_negedge_reg_1_sqmuxa_6_2,
       N_529,
       N_425,
       N_423,
       N_513,
       N_411,
       N_660,
       N_705,
       N_706,
       N_708,
       N_709,
       N_711,
       N_710,
       N_707,
       N_704,
       CoreAPB3_0_APBmslave0_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE,
       PRDATA_regif_sn_N_20_i_1,
       N_506,
       N_140,
       N_700,
       N_702,
       N_703,
       N_699,
       N_698
    );
input  [15:0] CoreAPB3_0_APBmslave0_PWDATA;
output [8:1] pwm_enable_reg;
output [128:1] pwm_negedge_reg;
output [15:0] period_reg;
input  [15:0] period_cnt;
output [5:5] PRDATA_regif_0_0;
input  [7:2] CoreAPB3_0_APBmslave0_PADDR;
output [1:1] PRDATA_regif_12_0;
output [4:4] PRDATA_regif_9_i_1;
output PRDATA_regif_9_i_0_4;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output N_428;
output N_629;
output N_678;
output N_689;
output N_686;
output N_679;
output N_687;
output N_688;
output N_690;
output N_680;
output N_685;
output N_681;
output N_684;
output N_691;
output psh_enable_reg1_1_sqmuxa_0;
output N_528;
output psh_negedge_reg_1_sqmuxa_6_2;
output N_529;
input  N_425;
input  N_423;
output N_513;
output N_411;
output N_660;
output N_705;
output N_706;
output N_708;
output N_709;
output N_711;
output N_710;
output N_707;
output N_704;
input  CoreAPB3_0_APBmslave0_PSELx;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;
output PRDATA_regif_sn_N_20_i_1;
output N_506;
output N_140;
output N_700;
output N_702;
output N_703;
output N_699;
output N_698;

    wire un1_period_cnt, un1_period_cnt_i_0, VCC_net_1, 
        psh_negedge_reg_1_sqmuxa_3_net_1, GND_net_1, 
        psh_negedge_reg_1_sqmuxa_2_net_1, 
        psh_negedge_reg_1_sqmuxa_1_net_1, 
        psh_negedge_reg_1_sqmuxa_net_1, psh_enable_reg1_1_sqmuxa, 
        psh_negedge_reg_1_sqmuxa_7_net_1, 
        psh_negedge_reg_1_sqmuxa_6_net_1, 
        psh_negedge_reg_1_sqmuxa_5_net_1, 
        psh_negedge_reg_1_sqmuxa_4_net_1, \psh_period_reg[3]_net_1 , 
        \psh_period_reg[4]_net_1 , \psh_period_reg[5]_net_1 , 
        \psh_period_reg[6]_net_1 , \psh_period_reg[7]_net_1 , 
        \psh_period_reg[8]_net_1 , \psh_period_reg[9]_net_1 , 
        \psh_period_reg[10]_net_1 , \psh_period_reg[11]_net_1 , 
        \psh_period_reg[12]_net_1 , \psh_period_reg[13]_net_1 , 
        \psh_period_reg[14]_net_1 , \psh_period_reg[15]_net_1 , 
        psh_period_reg_1_sqmuxa_net_1, \psh_period_reg[0]_net_1 , 
        \psh_period_reg[1]_net_1 , \psh_period_reg[2]_net_1 , 
        sync_update_net_1, sync_update_0_sqmuxa_net_1, 
        un1_period_cnt_cry_0, un1_period_cnt_cry_1, 
        un1_period_cnt_cry_2, un1_period_cnt_cry_3, 
        un1_period_cnt_cry_4, un1_period_cnt_cry_5, 
        un1_period_cnt_cry_6, un1_period_cnt_cry_7, 
        un1_period_cnt_cry_8, un1_period_cnt_cry_9, 
        un1_period_cnt_cry_10, un1_period_cnt_cry_11, 
        un1_period_cnt_cry_12, un1_period_cnt_cry_13, 
        un1_period_cnt_cry_14, N_433, \PRDATA_regif_0_0_1[5]_net_1 , 
        N_597, \PRDATA_regif_0_a2_1_0[5]_net_1 , N_431, N_659_1, 
        \PRDATA_regif_11_bm_1[0] , \PRDATA_regif_11_bm[0]_net_1 , 
        \PRDATA_regif_11_bm_1_1[11]_net_1 , 
        \PRDATA_regif_11_bm[11]_net_1 , 
        \PRDATA_regif_11_bm_1_1[8]_net_1 , 
        \PRDATA_regif_11_bm[8]_net_1 , \PRDATA_regif_11_bm_1[1] , 
        \PRDATA_regif_11_bm[1]_net_1 , 
        \PRDATA_regif_11_bm_1_1[9]_net_1 , 
        \PRDATA_regif_11_bm[9]_net_1 , 
        \PRDATA_regif_11_bm_1_1[10]_net_1 , 
        \PRDATA_regif_11_bm[10]_net_1 , \PRDATA_regif_11_am_1[2] , 
        \PRDATA_regif_11_am[2]_net_1 , \PRDATA_regif_11_bm_1[2] , 
        \PRDATA_regif_11_bm[2]_net_1 , \PRDATA_regif_11_am_1[7] , 
        \PRDATA_regif_11_am[7]_net_1 , \PRDATA_regif_11_bm_1[7] , 
        \PRDATA_regif_11_bm[7]_net_1 , \PRDATA_regif_11_am_1[3] , 
        \PRDATA_regif_11_am[3]_net_1 , \PRDATA_regif_11_bm_1[3] , 
        \PRDATA_regif_11_bm[3]_net_1 , \PRDATA_regif_11_am_1[6] , 
        \PRDATA_regif_11_am[6]_net_1 , \PRDATA_regif_11_bm_1[6] , 
        \PRDATA_regif_11_bm[6]_net_1 , 
        \PRDATA_regif_11_am_1_1[13]_net_1 , 
        \PRDATA_regif_11_am[13]_net_1 , 
        \PRDATA_regif_11_bm_1_1[13]_net_1 , 
        \PRDATA_regif_11_bm[13]_net_1 , \PRDATA_regif_0_m2_1_1[5] , 
        \PRDATA_regif_7_1[4] , \PRDATA_regif_11_am[0]_net_1 , 
        \PRDATA_regif_11_am[11]_net_1 , \PRDATA_regif_11_am[8]_net_1 , 
        \PRDATA_regif_11_am[1]_net_1 , \PRDATA_regif_11_am[9]_net_1 , 
        \PRDATA_regif_11_am[10]_net_1 , \PRDATA_regif_11_bm[12]_net_1 , 
        \PRDATA_regif_11_am[12]_net_1 , psh_period_reg_1_sqmuxa_2_0, 
        psh_negedge_reg_1_sqmuxa_2_0_0_net_1, 
        psh_negedge_reg_1_sqmuxa_1_0_0_net_1, 
        psh_negedge_reg_1_sqmuxa_0_net_1, N_424, N_611, N_612, N_613, 
        N_615, N_616, N_586, N_598, psh_negedge_reg_1_sqmuxa_7_1_net_1, 
        psh_negedge_reg_1_sqmuxa_3_1_net_1, 
        sync_update_0_sqmuxa_0_net_1, N_401, N_649, N_638, N_366, 
        N_629_0, N_625, N_646, N_644, N_672, N_654, N_653, N_634, 
        N_633, N_368, N_632, N_404, N_655, 
        \PRDATA_regif_9_i_0[0]_net_1 , \PRDATA_regif_9_i_0[12]_net_1 , 
        \PRDATA_regif_9_i_0[1]_net_1 , 
        \PRDATA_regif_9_i_m2_i_0[9]_net_1 , 
        \PRDATA_regif_9_i_0[10]_net_1 , \PRDATA_regif_9_i_0[8]_net_1 , 
        \PRDATA_regif_9_i_0[11]_net_1 , \PRDATA_regif_7_i_0[12]_net_1 , 
        psh_prescale_reg13_net_1;
    
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[70]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[70]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[42]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[42]));
    SLE \period_reg[5]  (.D(\psh_period_reg[5]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[5]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[27]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[27]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[126]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[126]));
    SLE \period_reg[14]  (.D(\psh_period_reg[14]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[14]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[111]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[111]));
    CFG2 #( .INIT(4'h8) )  psh_negedge_reg_1_sqmuxa_6_2_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        psh_negedge_reg_1_sqmuxa_6_2));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_15  (.A(period_reg[15])
        , .B(period_cnt[15]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_14), .S(), .Y(), .FCO(un1_period_cnt));
    CFG4 #( .INIT(16'h503F) )  
        \gen_pos_neg_shregs[6].psh_negedge_reg_RNIBNPE1[85]  (.A(
        pwm_negedge_reg[85]), .B(pwm_negedge_reg[69]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_7_1[4] ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[45]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[45]));
    CFG2 #( .INIT(4'h2) )  psh_enable_reg1_1_sqmuxa_0_inst_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(psh_enable_reg1_1_sqmuxa_0)
        );
    SLE \period_reg[12]  (.D(\psh_period_reg[12]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[12]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_8  (.A(period_reg[8]), 
        .B(period_cnt[8]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_7), .S(), .Y(), .FCO(un1_period_cnt_cry_8));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[82]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[82]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[0]  (.A(
        pwm_negedge_reg[113]), .B(pwm_negedge_reg[17]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[0]_net_1 ));
    CFG4 #( .INIT(16'h3050) )  \PRDATA_regif_11_i_a2[15]  (.A(
        pwm_negedge_reg[32]), .B(pwm_negedge_reg[96]), .C(
        psh_negedge_reg_1_sqmuxa_6_2), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_632));
    SLE \psh_period_reg[14]  (.D(CoreAPB3_0_APBmslave0_PWDATA[14]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[14]_net_1 )
        );
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[89]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[89]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[57]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[57]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[69]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[69]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[11]  (.A(
        pwm_negedge_reg[124]), .B(pwm_negedge_reg[28]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[11]_net_1 ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[1]  (.A(
        pwm_negedge_reg[50]), .B(pwm_negedge_reg[34]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[1] ));
    CFG4 #( .INIT(16'h1000) )  psh_negedge_reg_1_sqmuxa_3 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        psh_negedge_reg_1_sqmuxa_3_1_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_3_net_1)
        );
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[79]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[79]));
    SLE \period_reg[13]  (.D(\psh_period_reg[13]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[13]));
    CFG4 #( .INIT(16'h0020) )  psh_negedge_reg_1_sqmuxa_4 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_period_reg_1_sqmuxa_2_0), .D(N_528), .Y(
        psh_negedge_reg_1_sqmuxa_4_net_1));
    SLE \period_reg[8]  (.D(\psh_period_reg[8]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[8]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[101]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[101]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[20]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[20]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[7]  (.A(
        pwm_negedge_reg[56]), .B(pwm_negedge_reg[40]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[7] ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_am_1_1[7]  (.A(
        pwm_negedge_reg[120]), .B(pwm_negedge_reg[104]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_am_1[7] ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[3]  (.A(
        pwm_negedge_reg[52]), .B(pwm_negedge_reg[36]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[3] ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_am_1_1[3]  (.A(
        pwm_negedge_reg[116]), .B(pwm_negedge_reg[100]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_am_1[3] ));
    SLE \period_reg[11]  (.D(\psh_period_reg[11]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[11]));
    SLE \psh_period_reg[12]  (.D(CoreAPB3_0_APBmslave0_PWDATA[12]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[12]_net_1 )
        );
    SLE \psh_enable_reg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[4]));
    CFG4 #( .INIT(16'h3050) )  \PRDATA_regif_11_i_a2[14]  (.A(
        pwm_negedge_reg[31]), .B(pwm_negedge_reg[95]), .C(
        psh_negedge_reg_1_sqmuxa_6_2), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_653));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[92]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[92]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[97]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[97]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[37]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[37]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[8]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[8]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[23]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[23]));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_am[9]  (.A(N_638), .B(
        pwm_negedge_reg[10]), .C(\PRDATA_regif_9_i_m2_i_0[9]_net_1 ), 
        .D(N_425), .Y(\PRDATA_regif_11_am[9]_net_1 ));
    SLE \period_reg[3]  (.D(\psh_period_reg[3]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[3]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[65]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[65]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[119]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[119]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[105]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[105]));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_6[6]  (.A(pwm_enable_reg[7]), 
        .B(period_reg[6]), .C(CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        N_615));
    CFG4 #( .INIT(16'hC800) )  \PRDATA_regif_12[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_615), .C(N_431), .D(
        PRDATA_regif_sn_N_20_i_1), .Y(N_702));
    CFG4 #( .INIT(16'h8000) )  sync_update_0_sqmuxa_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        sync_update_0_sqmuxa_0_net_1));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[1]  (.A(
        pwm_negedge_reg[66]), .B(pwm_negedge_reg[82]), .C(
        \PRDATA_regif_11_bm_1[1] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[1]_net_1 ));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[46]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[46]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[9]  (.A(
        pwm_negedge_reg[58]), .B(pwm_negedge_reg[42]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_bm_1_1[9]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[75]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[75]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[11]  (.A(
        pwm_negedge_reg[60]), .B(pwm_negedge_reg[44]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_bm_1_1[11]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[2]  (.A(
        pwm_negedge_reg[67]), .B(pwm_negedge_reg[83]), .C(
        \PRDATA_regif_11_bm_1[2] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[2]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \PRDATA_regif_0_a2_1_1[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[7]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_659_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_14  (.A(period_reg[14])
        , .B(period_cnt[14]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_13), .S(), .Y(), .FCO(un1_period_cnt_cry_14)
        );
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[106]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[106]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[35]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[35]));
    SLE \psh_period_reg[8]  (.D(CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[8]_net_1 ));
    SLE \period_reg[0]  (.D(\psh_period_reg[0]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[0]));
    CFG4 #( .INIT(16'h0FAC) )  
        \gen_pos_neg_shregs[4].psh_negedge_reg_RNI32PC2[53]  (.A(
        pwm_negedge_reg[37]), .B(pwm_negedge_reg[53]), .C(
        \PRDATA_regif_7_1[4] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        N_629));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[0]_net_1 ), .C(
        \PRDATA_regif_11_am[0]_net_1 ), .Y(N_678));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[14]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[14]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_710));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[58]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[58]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[0]  (.A(
        pwm_negedge_reg[49]), .B(pwm_negedge_reg[33]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[0] ));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[10]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[10]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_706));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[7]  (.A(
        pwm_negedge_reg[72]), .B(pwm_negedge_reg[88]), .C(
        \PRDATA_regif_11_bm_1[7] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[7]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[114]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[114]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[60]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[60]));
    CFG4 #( .INIT(16'h0035) )  \PRDATA_regif_9_i_1[4]  (.A(
        pwm_negedge_reg[101]), .B(pwm_negedge_reg[5]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(PRDATA_regif_9_i_1[4]));
    CFG4 #( .INIT(16'h5030) )  \PRDATA_regif_11_i_a2_2[15]  (.A(
        pwm_negedge_reg[48]), .B(pwm_negedge_reg[112]), .C(N_423), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_634));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[44]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[44]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_1  (.A(period_reg[1]), 
        .B(period_cnt[1]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_0), .S(), .Y(), .FCO(un1_period_cnt_cry_1));
    CFG2 #( .INIT(4'h7) )  PRDATA_regif_sn_N_20_i_0_o2 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_528));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_am[0]  (.A(N_644), .B(
        pwm_negedge_reg[1]), .C(\PRDATA_regif_9_i_0[0]_net_1 ), .D(
        N_425), .Y(\PRDATA_regif_11_am[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_15_RNIHOI2  (.A(
        un1_period_cnt), .Y(un1_period_cnt_i_0));
    CFG2 #( .INIT(4'h8) )  psh_negedge_reg_1_sqmuxa_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        psh_negedge_reg_1_sqmuxa_0_net_1));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[118]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[118]));
    CFG4 #( .INIT(16'h0001) )  PRDATA_regif_sn_N_20_i_0_a2_3 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(N_672));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[87]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[87]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_11  (.A(period_reg[11])
        , .B(period_cnt[11]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_10), .S(), .Y(), .FCO(un1_period_cnt_cry_11)
        );
    SLE \psh_period_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[2]_net_1 ));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[80]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[80]));
    CFG4 #( .INIT(16'h1000) )  psh_enable_reg1_1_sqmuxa_2_0_RNI7NM71 (
        .A(CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_period_reg_1_sqmuxa_2_0), .D(psh_enable_reg1_1_sqmuxa_0), 
        .Y(psh_enable_reg1_1_sqmuxa));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[13]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[13]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_709));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[68]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[68]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[62]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[62]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[10]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[10]));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_bm[12]  (.A(N_625), .B(
        pwm_negedge_reg[77]), .C(\PRDATA_regif_7_i_0[12]_net_1 ), .D(
        N_425), .Y(\PRDATA_regif_11_bm[12]_net_1 ));
    CFG4 #( .INIT(16'h3050) )  \PRDATA_regif_11_i_a2_0[14]  (.A(
        pwm_negedge_reg[15]), .B(pwm_negedge_reg[79]), .C(N_425), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_654));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[78]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[78]));
    CFG2 #( .INIT(4'h8) )  psh_negedge_reg_1_sqmuxa_2_0_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        psh_negedge_reg_1_sqmuxa_2_0_0_net_1));
    SLE \psh_period_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[1]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_0_m2_0[5]  (.A(
        pwm_negedge_reg[22]), .B(pwm_negedge_reg[6]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_586));
    CFG4 #( .INIT(16'h503F) )  \PRDATA_regif_0_0_RNO_0[5]  (.A(
        pwm_negedge_reg[86]), .B(pwm_negedge_reg[70]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_0_m2_1_1[5] )
        );
    SLE \psh_period_reg[10]  (.D(CoreAPB3_0_APBmslave0_PWDATA[10]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[10]_net_1 )
        );
    CFG4 #( .INIT(16'hFFFE) )  \PRDATA_regif_11_i[15]  (.A(N_634), .B(
        N_633), .C(N_368), .D(N_632), .Y(N_506));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[8]  (.A(
        pwm_negedge_reg[73]), .B(pwm_negedge_reg[89]), .C(
        \PRDATA_regif_11_bm_1_1[8]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_bm[8]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[3]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[3]));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_am[13]  (.A(
        pwm_negedge_reg[14]), .B(pwm_negedge_reg[30]), .C(
        \PRDATA_regif_11_am_1_1[13]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_am[13]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_6[3]  (.A(pwm_enable_reg[4]), 
        .B(period_reg[3]), .C(CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        N_612));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[127]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[127]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[28]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[28]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[36]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[36]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_7  (.A(period_reg[7]), 
        .B(period_cnt[7]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_6), .S(), .Y(), .FCO(un1_period_cnt_cry_7));
    CFG3 #( .INIT(8'hE2) )  \PRDATA_regif_10_0_m2[0]  (.A(
        period_reg[0]), .B(CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        sync_update_net_1), .Y(N_598));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[22]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[22]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[10]  (.A(
        pwm_negedge_reg[123]), .B(pwm_negedge_reg[27]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[10]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[8]  (.A(
        pwm_negedge_reg[105]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_646));
    CFG3 #( .INIT(8'h80) )  sync_update_0_sqmuxa (.A(
        psh_prescale_reg13_net_1), .B(N_423), .C(
        sync_update_0_sqmuxa_0_net_1), .Y(sync_update_0_sqmuxa_net_1));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[10]  (.A(
        pwm_negedge_reg[59]), .B(pwm_negedge_reg[43]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_bm_1_1[10]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[11]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[11]_net_1 ), .C(
        \PRDATA_regif_11_am[11]_net_1 ), .Y(N_689));
    CFG4 #( .INIT(16'h5030) )  \PRDATA_regif_11_i_a2_1[15]  (.A(
        pwm_negedge_reg[64]), .B(pwm_negedge_reg[128]), .C(N_424), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_633));
    CFG4 #( .INIT(16'h0031) )  \PRDATA_regif_11_am[11]  (.A(N_425), .B(
        \PRDATA_regif_9_i_0[11]_net_1 ), .C(pwm_negedge_reg[12]), .D(
        N_401), .Y(\PRDATA_regif_11_am[11]_net_1 ));
    SLE \psh_period_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[0]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[15]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[15]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[84]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[84]));
    CFG4 #( .INIT(16'h0800) )  psh_negedge_reg_1_sqmuxa_3_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(
        CoreAPB3_0_APBmslave0_PADDR[7]), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(
        psh_negedge_reg_1_sqmuxa_3_1_net_1));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[4]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[4]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[34]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[34]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[11]  (.A(
        pwm_negedge_reg[108]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_401));
    CFG4 #( .INIT(16'hE4A0) )  \PRDATA_regif_10_0[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_598), .C(
        pwm_enable_reg[1]), .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(
        N_660));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[13]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[13]_net_1 ), .C(
        \PRDATA_regif_11_am[13]_net_1 ), .Y(N_691));
    SLE \period_reg[9]  (.D(\psh_period_reg[9]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[9]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[123]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[123]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[50]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[50]));
    SLE \period_reg[2]  (.D(\psh_period_reg[2]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[2]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_3  (.A(period_reg[3]), 
        .B(period_cnt[3]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_2), .S(), .Y(), .FCO(un1_period_cnt_cry_3));
    SLE \psh_period_reg[13]  (.D(CoreAPB3_0_APBmslave0_PWDATA[13]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[13]_net_1 )
        );
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[10]  (.A(
        pwm_negedge_reg[75]), .B(pwm_negedge_reg[91]), .C(
        \PRDATA_regif_11_bm_1_1[10]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_bm[10]_net_1 ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[94]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[94]));
    SLE \psh_enable_reg1[8]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[8]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[52]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[52]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[31]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[31]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[40]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[40]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[1]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[1]));
    CFG3 #( .INIT(8'hB8) )  \PRDATA_regif_11_ns[12]  (.A(
        \PRDATA_regif_11_bm[12]_net_1 ), .B(
        CoreAPB3_0_APBmslave0_PADDR[5]), .C(
        \PRDATA_regif_11_am[12]_net_1 ), .Y(N_690));
    SLE \psh_period_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[5]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[6]  (.A(
        pwm_negedge_reg[71]), .B(pwm_negedge_reg[87]), .C(
        \PRDATA_regif_11_bm_1[6] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[6]_net_1 ));
    CFG4 #( .INIT(16'hCCA0) )  \PRDATA_regif_12_0[1]  (.A(
        period_reg[1]), .B(pwm_enable_reg[2]), .C(N_431), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(PRDATA_regif_12_0[1]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_4  (.A(period_reg[4]), 
        .B(period_cnt[4]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_3), .S(), .Y(), .FCO(un1_period_cnt_cry_4));
    SLE sync_update (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(sync_update_0_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(sync_update_net_1));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_am[1]  (.A(N_629_0), 
        .B(pwm_negedge_reg[2]), .C(\PRDATA_regif_9_i_0[1]_net_1 ), .D(
        N_425), .Y(\PRDATA_regif_11_am[1]_net_1 ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[107]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[107]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[71]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[71]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[1]  (.A(
        pwm_negedge_reg[114]), .B(pwm_negedge_reg[18]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[1]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[3]  (.A(
        pwm_negedge_reg[68]), .B(pwm_negedge_reg[84]), .C(
        \PRDATA_regif_11_bm_1[3] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[3]_net_1 ));
    CFG4 #( .INIT(16'h0031) )  \PRDATA_regif_11_am[12]  (.A(N_425), .B(
        \PRDATA_regif_9_i_0[12]_net_1 ), .C(pwm_negedge_reg[13]), .D(
        N_366), .Y(\PRDATA_regif_11_am[12]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[7]_net_1 ), .C(
        \PRDATA_regif_11_am[7]_net_1 ), .Y(N_685));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_am[2]  (.A(
        pwm_negedge_reg[3]), .B(pwm_negedge_reg[19]), .C(
        \PRDATA_regif_11_am_1[2] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_am[2]_net_1 ));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_am[10]  (.A(N_649), .B(
        pwm_negedge_reg[11]), .C(\PRDATA_regif_9_i_0[10]_net_1 ), .D(
        N_425), .Y(\PRDATA_regif_11_am[10]_net_1 ));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[115]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[115]));
    CFG3 #( .INIT(8'h20) )  psh_negedge_reg_1_sqmuxa_7_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(N_431), .Y(
        psh_negedge_reg_1_sqmuxa_7_1_net_1));
    SLE \period_reg[4]  (.D(\psh_period_reg[4]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[4]));
    CFG4 #( .INIT(16'h8000) )  psh_negedge_reg_1_sqmuxa (.A(N_431), .B(
        psh_prescale_reg13_net_1), .C(N_659_1), .D(
        psh_negedge_reg_1_sqmuxa_0_net_1), .Y(
        psh_negedge_reg_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'hC800) )  \PRDATA_regif_12[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_613), .C(N_431), .D(
        PRDATA_regif_sn_N_20_i_1), .Y(N_700));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[116]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[116]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[43]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[43]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[13]  (.A(
        pwm_negedge_reg[62]), .B(pwm_negedge_reg[46]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_bm_1_1[13]_net_1 ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_am_1_1[13]  (.A(
        pwm_negedge_reg[126]), .B(pwm_negedge_reg[110]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_am_1_1[13]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  PRDATA_regif_sn_N_20_i_0 (.A(N_528), .B(
        N_423), .C(sync_update_0_sqmuxa_0_net_1), .D(N_672), .Y(
        PRDATA_regif_sn_N_20_i_1));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_am[7]  (.A(
        pwm_negedge_reg[8]), .B(pwm_negedge_reg[24]), .C(
        \PRDATA_regif_11_am_1[7] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_am[7]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[2]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[2]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[85]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[85]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[9]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[9]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_m2_i_0[9]  (.A(
        pwm_negedge_reg[122]), .B(pwm_negedge_reg[26]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_m2_i_0[9]_net_1 ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[103]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[103]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[63]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[63]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[13]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[13]));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[12]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[12]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_708));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[88]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[88]));
    CFG3 #( .INIT(8'h7F) )  \PRDATA_regif_0_0_1[5]  (.A(
        \PRDATA_regif_0_a2_1_0[5]_net_1 ), .B(N_431), .C(N_659_1), .Y(
        \PRDATA_regif_0_0_1[5]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[64]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[64]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[73]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[73]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[11]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[11]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[120]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[120]));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[1]  (.A(
        pwm_negedge_reg[98]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_629_0));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[99]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[99]));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[6]_net_1 ), .C(
        \PRDATA_regif_11_am[6]_net_1 ), .Y(N_684));
    CFG3 #( .INIT(8'h10) )  psh_enable_reg1_1_sqmuxa_2_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(psh_prescale_reg13_net_1), 
        .Y(psh_period_reg_1_sqmuxa_2_0));
    CFG4 #( .INIT(16'hC800) )  \PRDATA_regif_12[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_612), .C(N_431), .D(
        PRDATA_regif_sn_N_20_i_1), .Y(N_699));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[95]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[95]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_2  (.A(period_reg[2]), 
        .B(period_cnt[2]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_1), .S(), .Y(), .FCO(un1_period_cnt_cry_2));
    SLE \psh_period_reg[11]  (.D(CoreAPB3_0_APBmslave0_PWDATA[11]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[11]_net_1 )
        );
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[12]  (.A(
        pwm_negedge_reg[109]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_366));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[8]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[8]_net_1 ), .C(
        \PRDATA_regif_11_am[8]_net_1 ), .Y(N_686));
    CFG4 #( .INIT(16'h0405) )  \PRDATA_regif_11_am[8]  (.A(N_646), .B(
        pwm_negedge_reg[9]), .C(\PRDATA_regif_9_i_0[8]_net_1 ), .D(
        N_425), .Y(\PRDATA_regif_11_am[8]_net_1 ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[8]  (.A(
        pwm_negedge_reg[57]), .B(pwm_negedge_reg[41]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_11_bm_1_1[8]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_5  (.A(period_reg[5]), 
        .B(period_cnt[5]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_4), .S(), .Y(), .FCO(un1_period_cnt_cry_5));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[25]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[25]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[12]  (.A(
        pwm_negedge_reg[125]), .B(pwm_negedge_reg[29]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[12]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_12  (.A(period_reg[12])
        , .B(period_cnt[12]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_11), .S(), .Y(), .FCO(un1_period_cnt_cry_12)
        );
    CFG4 #( .INIT(16'hC0A0) )  \PRDATA_regif_0_a2_1_0[5]  (.A(
        pwm_negedge_reg[102]), .B(pwm_negedge_reg[118]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_0_a2_1_0[5]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \PRDATA_regif_0_a2_3[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(N_428));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[33]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[33]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[55]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[55]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[41]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[41]));
    CFG2 #( .INIT(4'h2) )  psh_negedge_reg_1_sqmuxa_1_0_0 (.A(
        CoreAPB3_0_APBmslave0_PADDR[6]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .Y(
        psh_negedge_reg_1_sqmuxa_1_0_0_net_1));
    CFG4 #( .INIT(16'h5030) )  \PRDATA_regif_11_i_a2_2[14]  (.A(
        pwm_negedge_reg[47]), .B(pwm_negedge_reg[111]), .C(N_423), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_655));
    CFG4 #( .INIT(16'hC800) )  \PRDATA_regif_12[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_616), .C(N_431), .D(
        PRDATA_regif_sn_N_20_i_1), .Y(N_703));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[19]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[19]));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[13]  (.A(
        pwm_negedge_reg[78]), .B(pwm_negedge_reg[94]), .C(
        \PRDATA_regif_11_bm_1_1[13]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_bm[13]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[49]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[49]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[110]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[110]));
    CFG4 #( .INIT(16'h8000) )  psh_negedge_reg_1_sqmuxa_6 (.A(N_428), 
        .B(psh_negedge_reg_1_sqmuxa_6_2), .C(psh_prescale_reg13_net_1), 
        .D(N_431), .Y(psh_negedge_reg_1_sqmuxa_6_net_1));
    SLE \psh_enable_reg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[7]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[122]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[122]));
    CFG4 #( .INIT(16'h0FAC) )  \PRDATA_regif_0_0_RNO[5]  (.A(
        pwm_negedge_reg[38]), .B(pwm_negedge_reg[54]), .C(
        \PRDATA_regif_0_m2_1_1[5] ), .D(CoreAPB3_0_APBmslave0_PADDR[4])
        , .Y(N_597));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[8]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[8]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_704));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[81]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[81]));
    SLE \psh_period_reg[9]  (.D(CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[9]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[15]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[15]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_711));
    CFG2 #( .INIT(4'hE) )  PRDATA_regif_sn_m23_i_o2 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_529));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[39]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[39]));
    SLE \period_reg[1]  (.D(\psh_period_reg[1]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[1]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[66]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[66]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_13  (.A(period_reg[13])
        , .B(period_cnt[13]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_12), .S(), .Y(), .FCO(un1_period_cnt_cry_13)
        );
    SLE \period_reg[6]  (.D(\psh_period_reg[6]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[6]));
    SLE \psh_enable_reg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[1]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[30]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[30]));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[9]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[9]_net_1 ), .C(
        \PRDATA_regif_11_am[9]_net_1 ), .Y(N_687));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[9]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[9]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_705));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[7]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[7]));
    CFG4 #( .INIT(16'h8000) )  psh_negedge_reg_1_sqmuxa_1 (.A(N_423), 
        .B(psh_negedge_reg_1_sqmuxa_1_0_0_net_1), .C(
        psh_prescale_reg13_net_1), .D(N_431), .Y(
        psh_negedge_reg_1_sqmuxa_1_net_1));
    CFG4 #( .INIT(16'hC800) )  \PRDATA_regif_12[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_611), .C(N_431), .D(
        PRDATA_regif_sn_N_20_i_1), .Y(N_698));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[76]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[76]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[17]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[17]));
    CFG2 #( .INIT(4'h8) )  PRDATA_regif_sn_N_20_i_0_a2_2 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_433));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[8]  (.A(
        pwm_negedge_reg[121]), .B(pwm_negedge_reg[25]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_9_i_0[8]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[53]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[53]));
    SLE \psh_enable_reg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[5]));
    SLE \psh_enable_reg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[3]));
    SLE \psh_enable_reg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[2]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[100]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[100]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[54]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[54]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_0  (.A(period_reg[0]), 
        .B(period_cnt[0]), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(un1_period_cnt_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_9  (.A(period_reg[9]), 
        .B(period_cnt[9]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_8), .S(), .Y(), .FCO(un1_period_cnt_cry_9));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[83]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[83]));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[91]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[91]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[124]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[124]));
    CFG4 #( .INIT(16'h5030) )  \PRDATA_regif_11_i_a2_1[14]  (.A(
        pwm_negedge_reg[63]), .B(pwm_negedge_reg[127]), .C(N_424), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_404));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_am[6]  (.A(
        pwm_negedge_reg[7]), .B(pwm_negedge_reg[23]), .C(
        \PRDATA_regif_11_am_1[6] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_am[6]_net_1 ));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[12]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[12]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[61]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[61]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[112]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[112]));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_am[3]  (.A(
        pwm_negedge_reg[4]), .B(pwm_negedge_reg[20]), .C(
        \PRDATA_regif_11_am_1[3] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_am[3]_net_1 ));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[90]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[90]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[128]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[128]));
    CFG4 #( .INIT(16'hFDDF) )  PRDATA_regif_sn_m23_i (.A(
        CoreAPB3_0_APBmslave0_PADDR[2]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        CoreAPB3_0_APBmslave0_PADDR[6]), .D(N_529), .Y(N_513));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[117]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[117]));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[3]_net_1 ), .C(
        \PRDATA_regif_11_am[3]_net_1 ), .Y(N_681));
    SLE \psh_period_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \PRDATA_regif_7_i_a2_3[12]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(N_424));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_10  (.A(period_reg[10])
        , .B(period_cnt[10]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_9), .S(), .Y(), .FCO(un1_period_cnt_cry_10));
    CFG4 #( .INIT(16'hFFFE) )  \PRDATA_regif_11_i[14]  (.A(N_653), .B(
        N_654), .C(N_404), .D(N_655), .Y(N_140));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[93]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[93]));
    SLE \psh_period_reg[15]  (.D(CoreAPB3_0_APBmslave0_PWDATA[15]), 
        .CLK(GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[15]_net_1 )
        );
    CFG2 #( .INIT(4'h4) )  psh_period_reg_1_sqmuxa_1 (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_431));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[11]  (.A(
        pwm_negedge_reg[76]), .B(pwm_negedge_reg[92]), .C(
        \PRDATA_regif_11_bm_1_1[11]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_bm[11]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_6[4]  (.A(pwm_enable_reg[5]), 
        .B(period_reg[4]), .C(CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        N_613));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[102]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[102]));
    CFG4 #( .INIT(16'h5300) )  \PRDATA_regif_7_i_0[12]  (.A(
        pwm_negedge_reg[93]), .B(pwm_negedge_reg[61]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        \PRDATA_regif_7_i_0[12]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  psh_negedge_reg_1_sqmuxa_5 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_period_reg_1_sqmuxa_2_0), .D(N_433), .Y(
        psh_negedge_reg_1_sqmuxa_5_net_1));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[86]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[86]));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[1]_net_1 ), .C(
        \PRDATA_regif_11_am[1]_net_1 ), .Y(N_679));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[10]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[10]_net_1 ), .C(
        \PRDATA_regif_11_am[10]_net_1 ), .Y(N_688));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[21]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[21]));
    CFG4 #( .INIT(16'h3050) )  \PRDATA_regif_11_i_a2_0[15]  (.A(
        pwm_negedge_reg[16]), .B(pwm_negedge_reg[80]), .C(N_425), .D(
        CoreAPB3_0_APBmslave0_PADDR[5]), .Y(N_368));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[6]  (.A(
        pwm_negedge_reg[55]), .B(pwm_negedge_reg[39]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[6] ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_am_1_1[6]  (.A(
        pwm_negedge_reg[119]), .B(pwm_negedge_reg[103]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_am_1[6] ));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[113]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[113]));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[109]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[109]));
    CFG3 #( .INIT(8'h80) )  psh_prescale_reg13 (.A(
        CoreAPB3_0_APBmslave0_PSELx), .B(CoreAPB3_0_APBmslave0_PWRITE), 
        .C(CoreAPB3_0_APBmslave0_PENABLE), .Y(psh_prescale_reg13_net_1)
        );
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_6[7]  (.A(pwm_enable_reg[8]), 
        .B(period_reg[7]), .C(CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        N_616));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[9]  (.A(
        pwm_negedge_reg[74]), .B(pwm_negedge_reg[90]), .C(
        \PRDATA_regif_11_bm_1_1[9]_net_1 ), .D(
        CoreAPB3_0_APBmslave0_PADDR[4]), .Y(
        \PRDATA_regif_11_bm[9]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_regif_0_a2_0[5]  (.A(N_428), .B(
        N_431), .C(CoreAPB3_0_APBmslave0_PADDR[4]), .D(N_586), .Y(
        N_411));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[5]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[5]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[16]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[16]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[72]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[72]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[48]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[48]));
    ARI1 #( .INIT(20'h5AA55) )  
        \gen_pos_neg_regs[1].un1_period_cnt_cry_6  (.A(period_reg[6]), 
        .B(period_cnt[6]), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_period_cnt_cry_5), .S(), .Y(), .FCO(un1_period_cnt_cry_6));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[98]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[98]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[24]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[24]));
    SLE \psh_period_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[4]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_m2_i_a2_2[9]  (.A(
        pwm_negedge_reg[106]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_638));
    CFG3 #( .INIT(8'hAC) )  \PRDATA_regif_6[2]  (.A(pwm_enable_reg[3]), 
        .B(period_reg[2]), .C(CoreAPB3_0_APBmslave0_PADDR[3]), .Y(
        N_611));
    SLE \gen_pos_neg_shregs[6].psh_negedge_reg[96]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_2_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[96]));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_bm_1_1[2]  (.A(
        pwm_negedge_reg[51]), .B(pwm_negedge_reg[35]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_bm_1[2] ));
    CFG4 #( .INIT(16'h05F3) )  \PRDATA_regif_11_am_1_1[2]  (.A(
        pwm_negedge_reg[115]), .B(pwm_negedge_reg[99]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(\PRDATA_regif_11_am_1[2] ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[104]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[104]));
    CFG4 #( .INIT(16'h0080) )  psh_negedge_reg_1_sqmuxa_2 (.A(N_428), 
        .B(psh_prescale_reg13_net_1), .C(
        psh_negedge_reg_1_sqmuxa_2_0_0_net_1), .D(N_528), .Y(
        psh_negedge_reg_1_sqmuxa_2_net_1));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[32]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[15]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[32]));
    CFG4 #( .INIT(16'h1000) )  psh_negedge_reg_1_sqmuxa_7 (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[6]), .C(
        psh_negedge_reg_1_sqmuxa_7_1_net_1), .D(
        psh_prescale_reg13_net_1), .Y(psh_negedge_reg_1_sqmuxa_7_net_1)
        );
    SLE \period_reg[7]  (.D(\psh_period_reg[7]_net_1 ), .CLK(GL0_INST), 
        .EN(un1_period_cnt_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(period_reg[7]));
    CFG4 #( .INIT(16'h3500) )  \PRDATA_regif_9_i_0[4]  (.A(
        pwm_negedge_reg[117]), .B(pwm_negedge_reg[21]), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(PRDATA_regif_9_i_0_4));
    SLE \psh_period_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[7]_net_1 ));
    SLE \gen_pos_neg_shregs[7].psh_negedge_reg[108]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[11]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_1_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[108]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[74]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[74]));
    CFG4 #( .INIT(16'hAC0F) )  \PRDATA_regif_11_bm[0]  (.A(
        pwm_negedge_reg[65]), .B(pwm_negedge_reg[81]), .C(
        \PRDATA_regif_11_bm_1[0] ), .D(CoreAPB3_0_APBmslave0_PADDR[4]), 
        .Y(\PRDATA_regif_11_bm[0]_net_1 ));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[51]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[51]));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[67]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[67]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[56]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[56]));
    SLE \period_reg[10]  (.D(\psh_period_reg[10]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[10]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[121]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[8]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[121]));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_7_i_a2_2[12]  (.A(
        pwm_negedge_reg[45]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_625));
    SLE \gen_pos_neg_shregs[5].psh_negedge_reg[77]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_3_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[77]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[26]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[9]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[26]));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[29]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[29]));
    SLE \gen_pos_neg_shregs[4].psh_negedge_reg[59]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[10]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_4_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[59]));
    SLE \psh_enable_reg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), 
        .CLK(GL0_INST), .EN(psh_enable_reg1_1_sqmuxa), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_enable_reg[6]));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[10]  (.A(
        pwm_negedge_reg[107]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_649));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[6]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[6]));
    CFG4 #( .INIT(16'h8F0F) )  \PRDATA_regif_0_0[5]  (.A(N_433), .B(
        N_428), .C(\PRDATA_regif_0_0_1[5]_net_1 ), .D(N_597), .Y(
        PRDATA_regif_0_0[5]));
    SLE \gen_pos_neg_shregs[1].psh_negedge_reg[14]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[13]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_7_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[14]));
    CFG4 #( .INIT(16'h1000) )  psh_period_reg_1_sqmuxa (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(
        CoreAPB3_0_APBmslave0_PADDR[7]), .C(
        psh_period_reg_1_sqmuxa_2_0), .D(N_431), .Y(
        psh_period_reg_1_sqmuxa_net_1));
    SLE \psh_period_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(psh_period_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\psh_period_reg[6]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_regif_12[11]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(N_672), .C(period_reg[11]), 
        .D(CoreAPB3_0_APBmslave0_PADDR[2]), .Y(N_707));
    SLE \gen_pos_neg_shregs[2].psh_negedge_reg[18]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_6_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[18]));
    CFG3 #( .INIT(8'hD8) )  \PRDATA_regif_11_ns[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[5]), .B(
        \PRDATA_regif_11_bm[2]_net_1 ), .C(
        \PRDATA_regif_11_am[2]_net_1 ), .Y(N_680));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[47]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[14]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[47]));
    SLE \gen_pos_neg_shregs[8].psh_negedge_reg[125]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[12]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[125]));
    SLE \period_reg[15]  (.D(\psh_period_reg[15]_net_1 ), .CLK(
        GL0_INST), .EN(un1_period_cnt_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(period_reg[15]));
    SLE \gen_pos_neg_shregs[3].psh_negedge_reg[38]  (.D(
        CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(GL0_INST), .EN(
        psh_negedge_reg_1_sqmuxa_5_net_1), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(pwm_negedge_reg[38]));
    CFG3 #( .INIT(8'h01) )  \PRDATA_regif_9_i_a2_2[0]  (.A(
        pwm_negedge_reg[97]), .B(CoreAPB3_0_APBmslave0_PADDR[4]), .C(
        CoreAPB3_0_APBmslave0_PADDR[3]), .Y(N_644));
    
endmodule


module corepwm_Z4_layer0(
       CoreAPB3_0_APBmslave0_PWDATA,
       PRDATA_regif_0_0,
       CoreAPB3_0_APBmslave0_PADDR,
       PRDATA_regif_12_0,
       PRDATA_regif_9_i_1,
       PRDATA_regif_9_i_0,
       PWM_c,
       pwm_enable_reg_5,
       period_reg_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_428,
       N_629,
       N_678,
       N_689,
       N_686,
       N_679,
       N_687,
       N_688,
       N_690,
       N_680,
       N_685,
       N_681,
       N_684,
       N_691,
       psh_enable_reg1_1_sqmuxa_0,
       N_528,
       psh_negedge_reg_1_sqmuxa_6_2,
       N_529,
       N_425,
       N_423,
       N_513,
       N_411,
       N_660,
       N_705,
       N_706,
       N_708,
       N_709,
       N_711,
       N_710,
       N_707,
       N_704,
       CoreAPB3_0_APBmslave0_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE,
       PRDATA_regif_sn_N_20_i_1,
       N_506,
       N_140,
       N_700,
       N_702,
       N_703,
       N_699,
       N_698
    );
input  [15:0] CoreAPB3_0_APBmslave0_PWDATA;
output [5:5] PRDATA_regif_0_0;
input  [7:2] CoreAPB3_0_APBmslave0_PADDR;
output [1:1] PRDATA_regif_12_0;
output [4:4] PRDATA_regif_9_i_1;
output [4:4] PRDATA_regif_9_i_0;
output [8:1] PWM_c;
output pwm_enable_reg_5;
output period_reg_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output N_428;
output N_629;
output N_678;
output N_689;
output N_686;
output N_679;
output N_687;
output N_688;
output N_690;
output N_680;
output N_685;
output N_681;
output N_684;
output N_691;
output psh_enable_reg1_1_sqmuxa_0;
output N_528;
output psh_negedge_reg_1_sqmuxa_6_2;
output N_529;
input  N_425;
input  N_423;
output N_513;
output N_411;
output N_660;
output N_705;
output N_706;
output N_708;
output N_709;
output N_711;
output N_710;
output N_707;
output N_704;
input  CoreAPB3_0_APBmslave0_PSELx;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;
output PRDATA_regif_sn_N_20_i_1;
output N_506;
output N_140;
output N_700;
output N_702;
output N_703;
output N_699;
output N_698;

    wire \pwm_enable_reg[1] , \pwm_enable_reg[2] , \pwm_enable_reg[3] , 
        \pwm_enable_reg[4] , \pwm_enable_reg[5] , \pwm_enable_reg[7] , 
        \pwm_enable_reg[8] , \pwm_negedge_reg[1] , 
        \pwm_negedge_reg[2] , \pwm_negedge_reg[3] , 
        \pwm_negedge_reg[4] , \pwm_negedge_reg[5] , 
        \pwm_negedge_reg[6] , \pwm_negedge_reg[7] , 
        \pwm_negedge_reg[8] , \pwm_negedge_reg[9] , 
        \pwm_negedge_reg[10] , \pwm_negedge_reg[11] , 
        \pwm_negedge_reg[12] , \pwm_negedge_reg[13] , 
        \pwm_negedge_reg[14] , \pwm_negedge_reg[15] , 
        \pwm_negedge_reg[16] , \pwm_negedge_reg[17] , 
        \pwm_negedge_reg[18] , \pwm_negedge_reg[19] , 
        \pwm_negedge_reg[20] , \pwm_negedge_reg[21] , 
        \pwm_negedge_reg[22] , \pwm_negedge_reg[23] , 
        \pwm_negedge_reg[24] , \pwm_negedge_reg[25] , 
        \pwm_negedge_reg[26] , \pwm_negedge_reg[27] , 
        \pwm_negedge_reg[28] , \pwm_negedge_reg[29] , 
        \pwm_negedge_reg[30] , \pwm_negedge_reg[31] , 
        \pwm_negedge_reg[32] , \pwm_negedge_reg[33] , 
        \pwm_negedge_reg[34] , \pwm_negedge_reg[35] , 
        \pwm_negedge_reg[36] , \pwm_negedge_reg[37] , 
        \pwm_negedge_reg[38] , \pwm_negedge_reg[39] , 
        \pwm_negedge_reg[40] , \pwm_negedge_reg[41] , 
        \pwm_negedge_reg[42] , \pwm_negedge_reg[43] , 
        \pwm_negedge_reg[44] , \pwm_negedge_reg[45] , 
        \pwm_negedge_reg[46] , \pwm_negedge_reg[47] , 
        \pwm_negedge_reg[48] , \pwm_negedge_reg[49] , 
        \pwm_negedge_reg[50] , \pwm_negedge_reg[51] , 
        \pwm_negedge_reg[52] , \pwm_negedge_reg[53] , 
        \pwm_negedge_reg[54] , \pwm_negedge_reg[55] , 
        \pwm_negedge_reg[56] , \pwm_negedge_reg[57] , 
        \pwm_negedge_reg[58] , \pwm_negedge_reg[59] , 
        \pwm_negedge_reg[60] , \pwm_negedge_reg[61] , 
        \pwm_negedge_reg[62] , \pwm_negedge_reg[63] , 
        \pwm_negedge_reg[64] , \pwm_negedge_reg[65] , 
        \pwm_negedge_reg[66] , \pwm_negedge_reg[67] , 
        \pwm_negedge_reg[68] , \pwm_negedge_reg[69] , 
        \pwm_negedge_reg[70] , \pwm_negedge_reg[71] , 
        \pwm_negedge_reg[72] , \pwm_negedge_reg[73] , 
        \pwm_negedge_reg[74] , \pwm_negedge_reg[75] , 
        \pwm_negedge_reg[76] , \pwm_negedge_reg[77] , 
        \pwm_negedge_reg[78] , \pwm_negedge_reg[79] , 
        \pwm_negedge_reg[80] , \pwm_negedge_reg[81] , 
        \pwm_negedge_reg[82] , \pwm_negedge_reg[83] , 
        \pwm_negedge_reg[84] , \pwm_negedge_reg[85] , 
        \pwm_negedge_reg[86] , \pwm_negedge_reg[87] , 
        \pwm_negedge_reg[88] , \pwm_negedge_reg[89] , 
        \pwm_negedge_reg[90] , \pwm_negedge_reg[91] , 
        \pwm_negedge_reg[92] , \pwm_negedge_reg[93] , 
        \pwm_negedge_reg[94] , \pwm_negedge_reg[95] , 
        \pwm_negedge_reg[96] , \pwm_negedge_reg[97] , 
        \pwm_negedge_reg[98] , \pwm_negedge_reg[99] , 
        \pwm_negedge_reg[100] , \pwm_negedge_reg[101] , 
        \pwm_negedge_reg[102] , \pwm_negedge_reg[103] , 
        \pwm_negedge_reg[104] , \pwm_negedge_reg[105] , 
        \pwm_negedge_reg[106] , \pwm_negedge_reg[107] , 
        \pwm_negedge_reg[108] , \pwm_negedge_reg[109] , 
        \pwm_negedge_reg[110] , \pwm_negedge_reg[111] , 
        \pwm_negedge_reg[112] , \pwm_negedge_reg[113] , 
        \pwm_negedge_reg[114] , \pwm_negedge_reg[115] , 
        \pwm_negedge_reg[116] , \pwm_negedge_reg[117] , 
        \pwm_negedge_reg[118] , \pwm_negedge_reg[119] , 
        \pwm_negedge_reg[120] , \pwm_negedge_reg[121] , 
        \pwm_negedge_reg[122] , \pwm_negedge_reg[123] , 
        \pwm_negedge_reg[124] , \pwm_negedge_reg[125] , 
        \pwm_negedge_reg[126] , \pwm_negedge_reg[127] , 
        \pwm_negedge_reg[128] , \period_reg[0] , \period_reg[1] , 
        \period_reg[2] , \period_reg[3] , \period_reg[4] , 
        \period_reg[6] , \period_reg[7] , \period_reg[8] , 
        \period_reg[9] , \period_reg[10] , \period_reg[11] , 
        \period_reg[12] , \period_reg[13] , \period_reg[14] , 
        \period_reg[15] , \period_cnt[0] , \period_cnt[1] , 
        \period_cnt[2] , \period_cnt[3] , \period_cnt[4] , 
        \period_cnt[5] , \period_cnt[6] , \period_cnt[7] , 
        \period_cnt[8] , \period_cnt[9] , \period_cnt[10] , 
        \period_cnt[11] , \period_cnt[12] , \period_cnt[13] , 
        \period_cnt[14] , \period_cnt[15] , GND_net_1, VCC_net_1;
    
    pwm_gen_8s_16s_0 \genblk5.pwm_gen  (.PWM_c({PWM_c[8], PWM_c[7], 
        PWM_c[6], PWM_c[5], PWM_c[4], PWM_c[3], PWM_c[2], PWM_c[1]}), 
        .period_cnt({\period_cnt[15] , \period_cnt[14] , 
        \period_cnt[13] , \period_cnt[12] , \period_cnt[11] , 
        \period_cnt[10] , \period_cnt[9] , \period_cnt[8] , 
        \period_cnt[7] , \period_cnt[6] , \period_cnt[5] , 
        \period_cnt[4] , \period_cnt[3] , \period_cnt[2] , 
        \period_cnt[1] , \period_cnt[0] }), .pwm_negedge_reg({
        \pwm_negedge_reg[128] , \pwm_negedge_reg[127] , 
        \pwm_negedge_reg[126] , \pwm_negedge_reg[125] , 
        \pwm_negedge_reg[124] , \pwm_negedge_reg[123] , 
        \pwm_negedge_reg[122] , \pwm_negedge_reg[121] , 
        \pwm_negedge_reg[120] , \pwm_negedge_reg[119] , 
        \pwm_negedge_reg[118] , \pwm_negedge_reg[117] , 
        \pwm_negedge_reg[116] , \pwm_negedge_reg[115] , 
        \pwm_negedge_reg[114] , \pwm_negedge_reg[113] , 
        \pwm_negedge_reg[112] , \pwm_negedge_reg[111] , 
        \pwm_negedge_reg[110] , \pwm_negedge_reg[109] , 
        \pwm_negedge_reg[108] , \pwm_negedge_reg[107] , 
        \pwm_negedge_reg[106] , \pwm_negedge_reg[105] , 
        \pwm_negedge_reg[104] , \pwm_negedge_reg[103] , 
        \pwm_negedge_reg[102] , \pwm_negedge_reg[101] , 
        \pwm_negedge_reg[100] , \pwm_negedge_reg[99] , 
        \pwm_negedge_reg[98] , \pwm_negedge_reg[97] , 
        \pwm_negedge_reg[96] , \pwm_negedge_reg[95] , 
        \pwm_negedge_reg[94] , \pwm_negedge_reg[93] , 
        \pwm_negedge_reg[92] , \pwm_negedge_reg[91] , 
        \pwm_negedge_reg[90] , \pwm_negedge_reg[89] , 
        \pwm_negedge_reg[88] , \pwm_negedge_reg[87] , 
        \pwm_negedge_reg[86] , \pwm_negedge_reg[85] , 
        \pwm_negedge_reg[84] , \pwm_negedge_reg[83] , 
        \pwm_negedge_reg[82] , \pwm_negedge_reg[81] , 
        \pwm_negedge_reg[80] , \pwm_negedge_reg[79] , 
        \pwm_negedge_reg[78] , \pwm_negedge_reg[77] , 
        \pwm_negedge_reg[76] , \pwm_negedge_reg[75] , 
        \pwm_negedge_reg[74] , \pwm_negedge_reg[73] , 
        \pwm_negedge_reg[72] , \pwm_negedge_reg[71] , 
        \pwm_negedge_reg[70] , \pwm_negedge_reg[69] , 
        \pwm_negedge_reg[68] , \pwm_negedge_reg[67] , 
        \pwm_negedge_reg[66] , \pwm_negedge_reg[65] , 
        \pwm_negedge_reg[64] , \pwm_negedge_reg[63] , 
        \pwm_negedge_reg[62] , \pwm_negedge_reg[61] , 
        \pwm_negedge_reg[60] , \pwm_negedge_reg[59] , 
        \pwm_negedge_reg[58] , \pwm_negedge_reg[57] , 
        \pwm_negedge_reg[56] , \pwm_negedge_reg[55] , 
        \pwm_negedge_reg[54] , \pwm_negedge_reg[53] , 
        \pwm_negedge_reg[52] , \pwm_negedge_reg[51] , 
        \pwm_negedge_reg[50] , \pwm_negedge_reg[49] , 
        \pwm_negedge_reg[48] , \pwm_negedge_reg[47] , 
        \pwm_negedge_reg[46] , \pwm_negedge_reg[45] , 
        \pwm_negedge_reg[44] , \pwm_negedge_reg[43] , 
        \pwm_negedge_reg[42] , \pwm_negedge_reg[41] , 
        \pwm_negedge_reg[40] , \pwm_negedge_reg[39] , 
        \pwm_negedge_reg[38] , \pwm_negedge_reg[37] , 
        \pwm_negedge_reg[36] , \pwm_negedge_reg[35] , 
        \pwm_negedge_reg[34] , \pwm_negedge_reg[33] , 
        \pwm_negedge_reg[32] , \pwm_negedge_reg[31] , 
        \pwm_negedge_reg[30] , \pwm_negedge_reg[29] , 
        \pwm_negedge_reg[28] , \pwm_negedge_reg[27] , 
        \pwm_negedge_reg[26] , \pwm_negedge_reg[25] , 
        \pwm_negedge_reg[24] , \pwm_negedge_reg[23] , 
        \pwm_negedge_reg[22] , \pwm_negedge_reg[21] , 
        \pwm_negedge_reg[20] , \pwm_negedge_reg[19] , 
        \pwm_negedge_reg[18] , \pwm_negedge_reg[17] , 
        \pwm_negedge_reg[16] , \pwm_negedge_reg[15] , 
        \pwm_negedge_reg[14] , \pwm_negedge_reg[13] , 
        \pwm_negedge_reg[12] , \pwm_negedge_reg[11] , 
        \pwm_negedge_reg[10] , \pwm_negedge_reg[9] , 
        \pwm_negedge_reg[8] , \pwm_negedge_reg[7] , 
        \pwm_negedge_reg[6] , \pwm_negedge_reg[5] , 
        \pwm_negedge_reg[4] , \pwm_negedge_reg[3] , 
        \pwm_negedge_reg[2] , \pwm_negedge_reg[1] }), .pwm_enable_reg({
        \pwm_enable_reg[8] , \pwm_enable_reg[7] , pwm_enable_reg_5, 
        \pwm_enable_reg[5] , \pwm_enable_reg[4] , \pwm_enable_reg[3] , 
        \pwm_enable_reg[2] , \pwm_enable_reg[1] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    timebase_16s \genblk4.genblk1.timebase  (.period_cnt({
        \period_cnt[15] , \period_cnt[14] , \period_cnt[13] , 
        \period_cnt[12] , \period_cnt[11] , \period_cnt[10] , 
        \period_cnt[9] , \period_cnt[8] , \period_cnt[7] , 
        \period_cnt[6] , \period_cnt[5] , \period_cnt[4] , 
        \period_cnt[3] , \period_cnt[2] , \period_cnt[1] , 
        \period_cnt[0] }), .period_reg({\period_reg[15] , 
        \period_reg[14] , \period_reg[13] , \period_reg[12] , 
        \period_reg[11] , \period_reg[10] , \period_reg[9] , 
        \period_reg[8] , \period_reg[7] , \period_reg[6] , 
        period_reg_5, \period_reg[4] , \period_reg[3] , 
        \period_reg[2] , \period_reg[1] , \period_reg[0] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST));
    reg_if_Z5_layer0 \genblk2.reg_if  (.CoreAPB3_0_APBmslave0_PWDATA({
        CoreAPB3_0_APBmslave0_PWDATA[15], 
        CoreAPB3_0_APBmslave0_PWDATA[14], 
        CoreAPB3_0_APBmslave0_PWDATA[13], 
        CoreAPB3_0_APBmslave0_PWDATA[12], 
        CoreAPB3_0_APBmslave0_PWDATA[11], 
        CoreAPB3_0_APBmslave0_PWDATA[10], 
        CoreAPB3_0_APBmslave0_PWDATA[9], 
        CoreAPB3_0_APBmslave0_PWDATA[8], 
        CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .pwm_enable_reg({
        \pwm_enable_reg[8] , \pwm_enable_reg[7] , pwm_enable_reg_5, 
        \pwm_enable_reg[5] , \pwm_enable_reg[4] , \pwm_enable_reg[3] , 
        \pwm_enable_reg[2] , \pwm_enable_reg[1] }), .pwm_negedge_reg({
        \pwm_negedge_reg[128] , \pwm_negedge_reg[127] , 
        \pwm_negedge_reg[126] , \pwm_negedge_reg[125] , 
        \pwm_negedge_reg[124] , \pwm_negedge_reg[123] , 
        \pwm_negedge_reg[122] , \pwm_negedge_reg[121] , 
        \pwm_negedge_reg[120] , \pwm_negedge_reg[119] , 
        \pwm_negedge_reg[118] , \pwm_negedge_reg[117] , 
        \pwm_negedge_reg[116] , \pwm_negedge_reg[115] , 
        \pwm_negedge_reg[114] , \pwm_negedge_reg[113] , 
        \pwm_negedge_reg[112] , \pwm_negedge_reg[111] , 
        \pwm_negedge_reg[110] , \pwm_negedge_reg[109] , 
        \pwm_negedge_reg[108] , \pwm_negedge_reg[107] , 
        \pwm_negedge_reg[106] , \pwm_negedge_reg[105] , 
        \pwm_negedge_reg[104] , \pwm_negedge_reg[103] , 
        \pwm_negedge_reg[102] , \pwm_negedge_reg[101] , 
        \pwm_negedge_reg[100] , \pwm_negedge_reg[99] , 
        \pwm_negedge_reg[98] , \pwm_negedge_reg[97] , 
        \pwm_negedge_reg[96] , \pwm_negedge_reg[95] , 
        \pwm_negedge_reg[94] , \pwm_negedge_reg[93] , 
        \pwm_negedge_reg[92] , \pwm_negedge_reg[91] , 
        \pwm_negedge_reg[90] , \pwm_negedge_reg[89] , 
        \pwm_negedge_reg[88] , \pwm_negedge_reg[87] , 
        \pwm_negedge_reg[86] , \pwm_negedge_reg[85] , 
        \pwm_negedge_reg[84] , \pwm_negedge_reg[83] , 
        \pwm_negedge_reg[82] , \pwm_negedge_reg[81] , 
        \pwm_negedge_reg[80] , \pwm_negedge_reg[79] , 
        \pwm_negedge_reg[78] , \pwm_negedge_reg[77] , 
        \pwm_negedge_reg[76] , \pwm_negedge_reg[75] , 
        \pwm_negedge_reg[74] , \pwm_negedge_reg[73] , 
        \pwm_negedge_reg[72] , \pwm_negedge_reg[71] , 
        \pwm_negedge_reg[70] , \pwm_negedge_reg[69] , 
        \pwm_negedge_reg[68] , \pwm_negedge_reg[67] , 
        \pwm_negedge_reg[66] , \pwm_negedge_reg[65] , 
        \pwm_negedge_reg[64] , \pwm_negedge_reg[63] , 
        \pwm_negedge_reg[62] , \pwm_negedge_reg[61] , 
        \pwm_negedge_reg[60] , \pwm_negedge_reg[59] , 
        \pwm_negedge_reg[58] , \pwm_negedge_reg[57] , 
        \pwm_negedge_reg[56] , \pwm_negedge_reg[55] , 
        \pwm_negedge_reg[54] , \pwm_negedge_reg[53] , 
        \pwm_negedge_reg[52] , \pwm_negedge_reg[51] , 
        \pwm_negedge_reg[50] , \pwm_negedge_reg[49] , 
        \pwm_negedge_reg[48] , \pwm_negedge_reg[47] , 
        \pwm_negedge_reg[46] , \pwm_negedge_reg[45] , 
        \pwm_negedge_reg[44] , \pwm_negedge_reg[43] , 
        \pwm_negedge_reg[42] , \pwm_negedge_reg[41] , 
        \pwm_negedge_reg[40] , \pwm_negedge_reg[39] , 
        \pwm_negedge_reg[38] , \pwm_negedge_reg[37] , 
        \pwm_negedge_reg[36] , \pwm_negedge_reg[35] , 
        \pwm_negedge_reg[34] , \pwm_negedge_reg[33] , 
        \pwm_negedge_reg[32] , \pwm_negedge_reg[31] , 
        \pwm_negedge_reg[30] , \pwm_negedge_reg[29] , 
        \pwm_negedge_reg[28] , \pwm_negedge_reg[27] , 
        \pwm_negedge_reg[26] , \pwm_negedge_reg[25] , 
        \pwm_negedge_reg[24] , \pwm_negedge_reg[23] , 
        \pwm_negedge_reg[22] , \pwm_negedge_reg[21] , 
        \pwm_negedge_reg[20] , \pwm_negedge_reg[19] , 
        \pwm_negedge_reg[18] , \pwm_negedge_reg[17] , 
        \pwm_negedge_reg[16] , \pwm_negedge_reg[15] , 
        \pwm_negedge_reg[14] , \pwm_negedge_reg[13] , 
        \pwm_negedge_reg[12] , \pwm_negedge_reg[11] , 
        \pwm_negedge_reg[10] , \pwm_negedge_reg[9] , 
        \pwm_negedge_reg[8] , \pwm_negedge_reg[7] , 
        \pwm_negedge_reg[6] , \pwm_negedge_reg[5] , 
        \pwm_negedge_reg[4] , \pwm_negedge_reg[3] , 
        \pwm_negedge_reg[2] , \pwm_negedge_reg[1] }), .period_reg({
        \period_reg[15] , \period_reg[14] , \period_reg[13] , 
        \period_reg[12] , \period_reg[11] , \period_reg[10] , 
        \period_reg[9] , \period_reg[8] , \period_reg[7] , 
        \period_reg[6] , period_reg_5, \period_reg[4] , 
        \period_reg[3] , \period_reg[2] , \period_reg[1] , 
        \period_reg[0] }), .period_cnt({\period_cnt[15] , 
        \period_cnt[14] , \period_cnt[13] , \period_cnt[12] , 
        \period_cnt[11] , \period_cnt[10] , \period_cnt[9] , 
        \period_cnt[8] , \period_cnt[7] , \period_cnt[6] , 
        \period_cnt[5] , \period_cnt[4] , \period_cnt[3] , 
        \period_cnt[2] , \period_cnt[1] , \period_cnt[0] }), 
        .PRDATA_regif_0_0({PRDATA_regif_0_0[5]}), 
        .CoreAPB3_0_APBmslave0_PADDR({CoreAPB3_0_APBmslave0_PADDR[7], 
        CoreAPB3_0_APBmslave0_PADDR[6], CoreAPB3_0_APBmslave0_PADDR[5], 
        CoreAPB3_0_APBmslave0_PADDR[4], CoreAPB3_0_APBmslave0_PADDR[3], 
        CoreAPB3_0_APBmslave0_PADDR[2]}), .PRDATA_regif_12_0({
        PRDATA_regif_12_0[1]}), .PRDATA_regif_9_i_1({
        PRDATA_regif_9_i_1[4]}), .PRDATA_regif_9_i_0_4(
        PRDATA_regif_9_i_0[4]), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .N_428(N_428)
        , .N_629(N_629), .N_678(N_678), .N_689(N_689), .N_686(N_686), 
        .N_679(N_679), .N_687(N_687), .N_688(N_688), .N_690(N_690), 
        .N_680(N_680), .N_685(N_685), .N_681(N_681), .N_684(N_684), 
        .N_691(N_691), .psh_enable_reg1_1_sqmuxa_0(
        psh_enable_reg1_1_sqmuxa_0), .N_528(N_528), 
        .psh_negedge_reg_1_sqmuxa_6_2(psh_negedge_reg_1_sqmuxa_6_2), 
        .N_529(N_529), .N_425(N_425), .N_423(N_423), .N_513(N_513), 
        .N_411(N_411), .N_660(N_660), .N_705(N_705), .N_706(N_706), 
        .N_708(N_708), .N_709(N_709), .N_711(N_711), .N_710(N_710), 
        .N_707(N_707), .N_704(N_704), .CoreAPB3_0_APBmslave0_PSELx(
        CoreAPB3_0_APBmslave0_PSELx), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .PRDATA_regif_sn_N_20_i_1(
        PRDATA_regif_sn_N_20_i_1), .N_506(N_506), .N_140(N_140), 
        .N_700(N_700), .N_702(N_702), .N_703(N_703), .N_699(N_699), 
        .N_698(N_698));
    
endmodule


module mss_sb_MSS(
       CoreAPB3_0_APBmslave0_PADDR,
       CoreAPB3_0_APBmslave0_PWDATA,
       COREI2C_0_0_INT,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_3,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_4,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_5,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_6,
       mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N,
       CoreAPB3_0_APBmslave0_PENABLE,
       mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave0_PWRITE,
       mss_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       CoreUARTapb_2_0_intr_or_2_Y,
       CoreUARTapb_2_1_intr_or_2_Y,
       CoreUARTapb_2_2_intr_or_2_Y,
       LOCK_0,
       GL0_INST
    );
output [8:0] CoreAPB3_0_APBmslave0_PADDR;
output [15:0] CoreAPB3_0_APBmslave0_PWDATA;
input  [0:0] COREI2C_0_0_INT;
input  [15:0] mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_3;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_4;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_5;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_6;
output mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N;
output CoreAPB3_0_APBmslave0_PENABLE;
output mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave0_PWRITE;
output mss_sb_MSS_TMP_0_MSS_RESET_N_M2F;
input  CoreUARTapb_2_0_intr_or_2_Y;
input  CoreUARTapb_2_1_intr_or_2_Y;
input  CoreUARTapb_2_2_intr_or_2_Y;
input  LOCK_0;
input  GL0_INST;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    MSS_010 #( .INIT(1438'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C00000000609300000003FFFFE400000000000010000000000F01C000001FEDFFC010842108421000001FE34001FF8000000400000000020051007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(0.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, 
        nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_6, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_5, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_4, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_3, nc56, nc57, nc58, 
        CoreAPB3_0_APBmslave0_PADDR[8], CoreAPB3_0_APBmslave0_PADDR[7], 
        CoreAPB3_0_APBmslave0_PADDR[6], CoreAPB3_0_APBmslave0_PADDR[5], 
        CoreAPB3_0_APBmslave0_PADDR[4], CoreAPB3_0_APBmslave0_PADDR[3], 
        CoreAPB3_0_APBmslave0_PADDR[2], CoreAPB3_0_APBmslave0_PADDR[1], 
        CoreAPB3_0_APBmslave0_PADDR[0]}), .F_HM0_ENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .F_HM0_SEL(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc59, 
        nc60}), .F_HM0_TRANS1(), .F_HM0_WDATA({nc61, nc62, nc63, nc64, 
        nc65, nc66, nc67, nc68, nc69, nc70, nc71, nc72, nc73, nc74, 
        nc75, nc76, CoreAPB3_0_APBmslave0_PWDATA[15], 
        CoreAPB3_0_APBmslave0_PWDATA[14], 
        CoreAPB3_0_APBmslave0_PWDATA[13], 
        CoreAPB3_0_APBmslave0_PWDATA[12], 
        CoreAPB3_0_APBmslave0_PWDATA[11], 
        CoreAPB3_0_APBmslave0_PWDATA[10], 
        CoreAPB3_0_APBmslave0_PWDATA[9], 
        CoreAPB3_0_APBmslave0_PWDATA[8], 
        CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc77, nc78}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc79, nc80, nc81, nc82}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc83, nc84}), .FAB_XDATAOUT({nc85, nc86, nc87, nc88, nc89, 
        nc90, nc91, nc92}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc93, 
        nc94}), .FIC32_1_MASTER({nc95, nc96}), .FPGA_RESET_N(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), .H2F_INTERRUPT({
        nc97, nc98, nc99, nc100, nc101, nc102, nc103, nc104, nc105, 
        nc106, nc107, nc108, nc109, nc110, nc111, nc112}), .H2F_NMI(), 
        .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc113, nc114, nc115, nc116, nc117, nc118, 
        nc119, nc120, nc121, nc122, nc123, nc124, nc125, nc126}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc127, nc128, nc129, nc130, nc131, nc132, 
        nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, nc141, 
        nc142, nc143, nc144, nc145, nc146, nc147, nc148, nc149, nc150, 
        nc151, nc152, nc153, nc154, nc155, nc156, nc157, nc158}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc159, nc160, nc161, nc162, 
        nc163, nc164, nc165, nc166, nc167, nc168}), .TRACECLK(), 
        .TRACEDATA({nc169, nc170, nc171, nc172}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc173, nc174, nc175, 
        nc176}), .TXDF({nc177, nc178, nc179, nc180, nc181, nc182, 
        nc183, nc184}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc185, nc186, nc187, nc188})
        , .F_BRESP_HRESP0({nc189, nc190}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc191, nc192, nc193, nc194, nc195, nc196, 
        nc197, nc198, nc199, nc200, nc201, nc202, nc203, nc204, nc205, 
        nc206, nc207, nc208, nc209, nc210, nc211, nc212, nc213, nc214, 
        nc215, nc216, nc217, nc218, nc219, nc220, nc221, nc222, nc223, 
        nc224, nc225, nc226, nc227, nc228, nc229, nc230, nc231, nc232, 
        nc233, nc234, nc235, nc236, nc237, nc238, nc239, nc240, nc241, 
        nc242, nc243, nc244, nc245, nc246, nc247, nc248, nc249, nc250, 
        nc251, nc252, nc253, nc254}), .F_RID({nc255, nc256, nc257, 
        nc258}), .F_RLAST(), .F_RRESP_HRESP1({nc259, nc260}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc261, nc262, 
        nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, nc271, 
        nc272, nc273, nc274, nc275, nc276}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        CoreUARTapb_2_2_intr_or_2_Y, CoreUARTapb_2_1_intr_or_2_Y, 
        CoreUARTapb_2_0_intr_or_2_Y, COREI2C_0_0_INT[0]}), .F2HCALIB(
        VCC_net_1), .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_FM0_ENABLE(GND_net_1), 
        .F_FM0_MASTLOCK(GND_net_1), .F_FM0_READY(VCC_net_1), 
        .F_FM0_SEL(GND_net_1), .F_FM0_SIZE({GND_net_1, GND_net_1}), 
        .F_FM0_TRANS1(GND_net_1), .F_FM0_WDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_FM0_WRITE(GND_net_1), .F_HM0_RDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1], 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0]}), .F_HM0_READY(
        VCC_net_1), .F_HM0_RESP(GND_net_1), .FAB_AVALID(VCC_net_1), 
        .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(LOCK_0), .FAB_RXACTIVE(VCC_net_1), 
        .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(GND_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(VCC_net_1), .XCLK_FAB(VCC_net_1), 
        .CLK_BASE(GL0_INST), .CLK_MDDR_APB(VCC_net_1), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), .SPI1_SCK_IN(
        GND_net_1), .SPI1_SDI_MGPIO11A_IN(GND_net_1), 
        .SPI1_SDO_MGPIO12A_IN(GND_net_1), .SPI1_SS0_MGPIO13A_IN(
        GND_net_1), .SPI1_SS1_MGPIO14A_IN(GND_net_1), 
        .SPI1_SS2_MGPIO15A_IN(GND_net_1), .SPI1_SS3_MGPIO16A_IN(
        GND_net_1), .SPI1_SS4_MGPIO17A_IN(GND_net_1), 
        .SPI1_SS5_MGPIO18A_IN(GND_net_1), .SPI1_SS6_MGPIO23A_IN(
        GND_net_1), .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc277, nc278, 
        nc279, nc280, nc281, nc282, nc283, nc284, nc285, nc286, nc287, 
        nc288, nc289, nc290, nc291, nc292}), .DRAM_BA({nc293, nc294, 
        nc295}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc296, nc297, nc298}), .DRAM_DQ_OUT({nc299, 
        nc300, nc301, nc302, nc303, nc304, nc305, nc306, nc307, nc308, 
        nc309, nc310, nc311, nc312, nc313, nc314, nc315, nc316}), 
        .DRAM_DQS_OUT({nc317, nc318, nc319}), .DRAM_FIFO_WE_OUT({nc320, 
        nc321}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc322, nc323, 
        nc324}), .DRAM_DQ_OE({nc325, nc326, nc327, nc328, nc329, nc330, 
        nc331, nc332, nc333, nc334, nc335, nc336, nc337, nc338, nc339, 
        nc340, nc341, nc342}), .DRAM_DQS_OE({nc343, nc344, nc345}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_2_Rx_async_1s_0s_1s_2s(
       rx_byte,
       controlReg2,
       clear_parity_reg,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       BT_TX_c,
       CoreUARTapb_2_2_PARITY_ERR,
       stop_strobe,
       CoreUARTapb_2_2_FRAMING_ERR,
       clear_parity_en,
       fifo_write,
       rx_idle
    );
output [7:0] rx_byte;
input  [2:0] controlReg2;
input  clear_parity_reg;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  baud_clock;
input  BT_TX_c;
output CoreUARTapb_2_2_PARITY_ERR;
output stop_strobe;
output CoreUARTapb_2_2_FRAMING_ERR;
output clear_parity_en;
output fifo_write;
output rx_idle;

    wire clear_parity_reg_i_0, \rx_bit_cnt[0]_net_1 , VCC_net_1, 
        \rx_bit_cnt_4[0] , GND_net_1, \rx_bit_cnt[1]_net_1 , 
        \rx_bit_cnt_4[1] , \rx_bit_cnt[2]_net_1 , \rx_bit_cnt_4[2] , 
        \rx_bit_cnt[3]_net_1 , \rx_bit_cnt_4[3] , \samples[1]_net_1 , 
        \samples[2]_net_1 , \rx_shift[0]_net_1 , \rx_shift_11[0] , 
        un1_samples7_1_0_2, \rx_shift[1]_net_1 , \rx_shift_11[1] , 
        \rx_shift[2]_net_1 , \rx_shift_11[2] , \rx_shift[3]_net_1 , 
        \rx_shift_11[3] , \rx_shift[4]_net_1 , \rx_shift_11[4] , 
        \rx_shift[5]_net_1 , \rx_shift_11[5] , \rx_shift[6]_net_1 , 
        \rx_shift_11[6] , \rx_shift[7]_net_1 , \rx_shift_11[7] , 
        \rx_shift[8]_net_1 , \rx_shift_11[8] , 
        \receive_count[0]_net_1 , N_373_i_0, \receive_count[1]_net_1 , 
        N_372_i_0, \receive_count[2]_net_1 , N_371_i_0, 
        \receive_count[3]_net_1 , N_370_i_0, clear_parity_en_9, 
        \rx_byte_2[7] , \samples[0]_net_1 , N_310, 
        parity_err_1_sqmuxa_i_0, rx_parity_calc_net_1, N_369_i_0, 
        framing_error_int_net_1, framing_error_int_0_sqmuxa, 
        framing_error_int_2_sqmuxa, framing_error_1_sqmuxa_i_0, 
        \rx_state[1]_net_1 , N_233_i_0, \rx_state[0]_net_1 , 
        \rx_state_ns[0] , clear_parity_en_9_i_0, rx_bit_cnt_1_sqmuxa, 
        rx_bit_cnt_0_sqmuxa, N_399, rx_state19_NE_1, N_243, 
        rx_state19_li, clear_parity_en_1_sqmuxa_net_1, 
        parity_err_0_sqmuxa_1_1_net_1, parity_err_0_sqmuxa_3_1_net_1, 
        clear_parity_en_0_sqmuxa_net_1, N_242, 
        framing_error_int_0_sqmuxa_0_a2_2_net_1, N_376, 
        framing_error_int5, N_403, parity_err_0_sqmuxa_1_net_1, 
        parity_err_0_sqmuxa_3_net_1, N_420, un1_parity_err31_1_net_1, 
        N_389, CO1;
    
    CFG4 #( .INIT(16'h4000) )  parity_err_0_sqmuxa_3 (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(
        parity_err_0_sqmuxa_3_1_net_1), .D(controlReg2[0]), .Y(
        parity_err_0_sqmuxa_3_net_1));
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[2]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  \rcv_cnt.receive_count_3_i_a2[0]  (.A(
        \receive_count[1]_net_1 ), .B(\receive_count[2]_net_1 ), .C(
        rx_idle), .D(\receive_count[3]_net_1 ), .Y(N_403));
    CFG3 #( .INIT(8'h20) )  framing_error_int_2_sqmuxa_0_a3 (.A(
        \receive_count[3]_net_1 ), .B(N_376), .C(\rx_state[1]_net_1 ), 
        .Y(framing_error_int_2_sqmuxa));
    CFG4 #( .INIT(16'hCCCE) )  un1_samples7_1_0 (.A(baud_clock), .B(
        rx_bit_cnt_1_sqmuxa), .C(\rx_state[0]_net_1 ), .D(
        \rx_state[1]_net_1 ), .Y(un1_samples7_1_0_2));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[0]));
    CFG4 #( .INIT(16'hE800) )  \rcv_cnt.receive_count_3_i_a2_0[3]  (.A(
        \samples[0]_net_1 ), .B(\samples[1]_net_1 ), .C(
        \samples[2]_net_1 ), .D(rx_idle), .Y(N_399));
    SLE \receive_count[1]  (.D(N_372_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[1]_net_1 ));
    SLE \rx_shift[7]  (.D(\rx_shift_11[7] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[7]_net_1 ));
    CFG4 #( .INIT(16'h1441) )  
        \make_parity_err.parity_err_12_iv_0_111_a2  (.A(
        clear_parity_reg), .B(framing_error_int5), .C(
        rx_parity_calc_net_1), .D(controlReg2[2]), .Y(N_310));
    CFG3 #( .INIT(8'h08) )  framing_error_int_0_sqmuxa_0_a2_2 (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(
        framing_error_int_0_sqmuxa_0_a2_2_net_1));
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  framing_error_RNO (.A(clear_parity_reg), .Y(
        clear_parity_reg_i_0));
    CFG2 #( .INIT(4'h8) )  clear_parity_en_0_sqmuxa (.A(controlReg2[0])
        , .B(controlReg2[1]), .Y(clear_parity_en_0_sqmuxa_net_1));
    CFG2 #( .INIT(4'h1) )  parity_err_0_sqmuxa_3_1 (.A(
        \rx_bit_cnt[1]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .Y(
        parity_err_0_sqmuxa_3_1_net_1));
    CFG3 #( .INIT(8'h10) )  rx_bit_cnt_0_sqmuxa_0_a3 (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .C(baud_clock), 
        .Y(rx_bit_cnt_0_sqmuxa));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[0]  (.A(rx_idle), 
        .B(\rx_shift[1]_net_1 ), .Y(\rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(N_370_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h1) )  \rx_state_ns_0_a3_0_3_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(\rx_state[0]_net_1 ), .Y(rx_idle));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[4]));
    CFG4 #( .INIT(16'hF7FF) )  un1_parity_err31_1 (.A(controlReg2[1]), 
        .B(\receive_count[3]_net_1 ), .C(N_376), .D(baud_clock), .Y(
        un1_parity_err31_1_net_1));
    CFG4 #( .INIT(16'h040E) )  \receive_shift.rx_shift_11[8]  (.A(
        clear_parity_en_0_sqmuxa_net_1), .B(\rx_shift[8]_net_1 ), .C(
        rx_idle), .D(framing_error_int5), .Y(\rx_shift_11[8] ));
    SLE rx_parity_calc (.D(N_369_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        rx_parity_calc_net_1));
    SLE \rx_bit_cnt[2]  (.D(\rx_bit_cnt_4[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[2]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[3]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(CO1), .D(
        rx_bit_cnt_0_sqmuxa), .Y(\rx_bit_cnt_4[3] ));
    SLE \rx_bit_cnt[1]  (.D(\rx_bit_cnt_4[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[1]_net_1 ));
    CFG3 #( .INIT(8'h21) )  rx_parity_calc_RNO (.A(
        rx_parity_calc_net_1), .B(\rx_state[1]_net_1 ), .C(N_389), .Y(
        N_369_i_0));
    CFG4 #( .INIT(16'h002E) )  \receive_shift.rx_shift_11[7]  (.A(
        N_242), .B(N_243), .C(framing_error_int5), .D(rx_idle), .Y(
        \rx_shift_11[7] ));
    CFG4 #( .INIT(16'h1230) )  \receive_count_RNO[2]  (.A(
        \receive_count[0]_net_1 ), .B(N_399), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_371_i_0));
    CFG3 #( .INIT(8'hAC) )  \receive_shift.rx_shift_9_0[7]  (.A(
        \rx_shift[8]_net_1 ), .B(\rx_shift[7]_net_1 ), .C(
        controlReg2[1]), .Y(N_242));
    CFG4 #( .INIT(16'h4002) )  \rcv_sm.rx_state19_NE_1  (.A(
        \rx_bit_cnt[3]_net_1 ), .B(\rx_bit_cnt[2]_net_1 ), .C(
        \rx_bit_cnt[1]_net_1 ), .D(clear_parity_en_1_sqmuxa_net_1), .Y(
        rx_state19_NE_1));
    SLE stop_strobe_inst_1 (.D(framing_error_int_2_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG4 #( .INIT(16'h0203) )  \rx_state_RNO[1]  (.A(
        \rx_state[1]_net_1 ), .B(rx_idle), .C(
        framing_error_int_2_sqmuxa), .D(rx_state19_li), .Y(N_233_i_0));
    CFG2 #( .INIT(4'h1) )  clear_parity_en_1_sqmuxa (.A(controlReg2[0])
        , .B(controlReg2[1]), .Y(clear_parity_en_1_sqmuxa_net_1));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[1]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[2]  (.A(rx_idle), 
        .B(\rx_shift[3]_net_1 ), .Y(\rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(N_371_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[2]_net_1 ));
    SLE clear_parity_en_1 (.D(clear_parity_en_9), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_en));
    CFG3 #( .INIT(8'h80) )  \un1_rx_bit_cnt_1.CO1  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_1_sqmuxa), .C(
        \rx_bit_cnt[1]_net_1 ), .Y(CO1));
    SLE \rx_state[1]  (.D(N_233_i_0), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[6]));
    CFG3 #( .INIT(8'h12) )  \receive_count_RNO[1]  (.A(
        \receive_count[0]_net_1 ), .B(N_399), .C(
        \receive_count[1]_net_1 ), .Y(N_372_i_0));
    GND GND (.Y(GND_net_1));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[3]  (.A(rx_idle), 
        .B(\rx_shift[4]_net_1 ), .Y(\rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(\rx_byte_2[7] ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[7]));
    CFG3 #( .INIT(8'hD7) )  \rcv_sm.rx_state19_NE  (.A(rx_state19_NE_1)
        , .B(\rx_bit_cnt[0]_net_1 ), .C(N_243), .Y(rx_state19_li));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[2]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(CO1), .Y(
        \rx_bit_cnt_4[2] ));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[3]));
    CFG3 #( .INIT(8'h40) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_0_a2  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9));
    CFG3 #( .INIT(8'h20) )  rx_bit_cnt_1_sqmuxa_0_a3 (.A(baud_clock), 
        .B(N_376), .C(\receive_count[3]_net_1 ), .Y(
        rx_bit_cnt_1_sqmuxa));
    CFG4 #( .INIT(16'h0009) )  \receive_count_RNO[3]  (.A(N_376), .B(
        \receive_count[3]_net_1 ), .C(N_399), .D(N_420), .Y(N_370_i_0));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[2]));
    CFG2 #( .INIT(4'h8) )  \rcv_sm.rx_byte_2[7]  (.A(controlReg2[0]), 
        .B(\rx_shift[7]_net_1 ), .Y(\rx_byte_2[7] ));
    CFG3 #( .INIT(8'h01) )  \receive_count_RNO[0]  (.A(N_399), .B(
        \receive_count[0]_net_1 ), .C(N_403), .Y(N_373_i_0));
    SLE parity_err (.D(N_310), .CLK(GL0_INST), .EN(
        parity_err_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_2_PARITY_ERR));
    SLE \rx_shift[6]  (.D(\rx_shift_11[6] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[6]_net_1 ));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[4]  (.A(rx_idle), 
        .B(\rx_shift[5]_net_1 ), .Y(\rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[3]_net_1 ));
    CFG4 #( .INIT(16'h040E) )  \receive_shift.rx_shift_11[6]  (.A(
        clear_parity_en_1_sqmuxa_net_1), .B(\rx_shift[7]_net_1 ), .C(
        rx_idle), .D(framing_error_int5), .Y(\rx_shift_11[6] ));
    CFG2 #( .INIT(4'h2) )  parity_err_0_sqmuxa_1_1 (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .Y(
        parity_err_0_sqmuxa_1_1_net_1));
    SLE framing_error_int (.D(framing_error_int_0_sqmuxa), .CLK(
        GL0_INST), .EN(baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(framing_error_int_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \rx_state_ns_0_0[0]  (.A(N_420), .B(
        rx_state19_li), .C(\rx_state[0]_net_1 ), .D(
        \receive_count[3]_net_1 ), .Y(\rx_state_ns[0] ));
    CFG4 #( .INIT(16'h0080) )  parity_err_0_sqmuxa_1 (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        parity_err_0_sqmuxa_1_1_net_1), .D(controlReg2[0]), .Y(
        parity_err_0_sqmuxa_1_net_1));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \samples[2]  (.D(BT_TX_c), .CLK(GL0_INST), .EN(baud_clock), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    SLE \receive_count[0]  (.D(N_373_i_0), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(GL0_INST), .EN(
        clear_parity_en_9), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_byte[5]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[5]  (.A(rx_idle), 
        .B(\rx_shift[6]_net_1 ), .Y(\rx_shift_11[5] ));
    CFG4 #( .INIT(16'h8000) )  framing_error_int_0_sqmuxa_0_a2 (.A(
        \receive_count[3]_net_1 ), .B(\rx_state[1]_net_1 ), .C(
        framing_error_int5), .D(
        framing_error_int_0_sqmuxa_0_a2_2_net_1), .Y(
        framing_error_int_0_sqmuxa));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[0]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(
        rx_bit_cnt_1_sqmuxa), .Y(\rx_bit_cnt_4[0] ));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[5]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \rcv_cnt.receive_count_3_i_o2[3]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(N_376));
    SLE \rx_bit_cnt[0]  (.D(\rx_bit_cnt_4[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[0]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  framing_error_1_sqmuxa_i (.A(
        framing_error_int_net_1), .B(clear_parity_reg), .C(baud_clock), 
        .Y(framing_error_1_sqmuxa_i_0));
    SLE \rx_shift[8]  (.D(\rx_shift_11[8] ), .CLK(GL0_INST), .EN(
        un1_samples7_1_0_2), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_shift[8]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[1]  (.A(rx_idle), 
        .B(\rx_shift[2]_net_1 ), .Y(\rx_shift_11[1] ));
    CFG3 #( .INIT(8'hBF) )  
        \receive_full_indicator.clear_parity_en_9_0_a3_0_a2_i  (.A(
        rx_state19_li), .B(\rx_state[0]_net_1 ), .C(baud_clock), .Y(
        clear_parity_en_9_i_0));
    CFG3 #( .INIT(8'h17) )  \rx_filtered.m3  (.A(\samples[1]_net_1 ), 
        .B(\samples[0]_net_1 ), .C(\samples[2]_net_1 ), .Y(
        framing_error_int5));
    SLE framing_error (.D(clear_parity_reg_i_0), .CLK(GL0_INST), .EN(
        framing_error_1_sqmuxa_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreUARTapb_2_2_FRAMING_ERR));
    CFG4 #( .INIT(16'hFFF7) )  \rx_par_calc.rx_parity_calc_4_u_i_o2  (
        .A(\receive_count[3]_net_1 ), .B(controlReg2[1]), .C(N_376), 
        .D(framing_error_int5), .Y(N_389));
    CFG2 #( .INIT(4'h6) )  \receive_shift.rx_shift_9_sn_m1  (.A(
        controlReg2[0]), .B(controlReg2[1]), .Y(N_243));
    CFG4 #( .INIT(16'h0004) )  \rcv_cnt.receive_count_3_i_a2_1[3]  (.A(
        \receive_count[0]_net_1 ), .B(rx_idle), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_420));
    CFG4 #( .INIT(16'hAAFE) )  parity_err_1_sqmuxa_i (.A(
        clear_parity_reg), .B(parity_err_0_sqmuxa_1_net_1), .C(
        parity_err_0_sqmuxa_3_net_1), .D(un1_parity_err31_1_net_1), .Y(
        parity_err_1_sqmuxa_i_0));
    SLE \rx_bit_cnt[3]  (.D(\rx_bit_cnt_4[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[1]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        rx_bit_cnt_1_sqmuxa), .D(rx_bit_cnt_0_sqmuxa), .Y(
        \rx_bit_cnt_4[1] ));
    
endmodule


module mss_sb_CoreUARTapb_2_2_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] tx_hold_reg;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, tx_hold_reg[7], 
        tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], tx_hold_reg[3], 
        tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]}), .C_WEN(
        INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), 
        .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({
        GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_2_fifo_ctrl_128(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_3636_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, \counter[0]_net_1 , 
        VCC_net_1, un1_counter_cry_0_Y_6, GND_net_1, 
        \counter[1]_net_1 , un1_counter_cry_1_0_S_5, 
        \counter[2]_net_1 , un1_counter_cry_2_0_S_5, 
        \counter[3]_net_1 , un1_counter_cry_3_0_S_5, 
        \counter[4]_net_1 , un1_counter_cry_4_0_S_5, 
        \counter[5]_net_1 , un1_counter_cry_5_0_S_5, 
        \counter[6]_net_1 , un1_counter_s_6_S_5, \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \data_out_0[0] , 
        \data_out_0[1] , \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_304_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_305_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        empty_4_net_1, full_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_305_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_2_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[2]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S_5), .Y(), .FCO(
        un1_counter_cry_2));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIJDO3 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_4_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[4]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S_5), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_304_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  full_4_RNIODH (.A(\counter[0]_net_1 ), 
        .B(full_4_net_1), .C(\counter[6]_net_1 ), .D(
        \counter[4]_net_1 ), .Y(fifo_full_tx_i_0));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[0]));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_305 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_305_FCO));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[6]));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_3_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[3]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S_5), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_tx), .C(fifo_write_tx), .D(
        GND_net_1), .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_6), 
        .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_3636_i_0 (.A(fifo_write_tx), .Y(
        N_3636_i_0_net_1));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[4]_net_1 ), 
        .Y(fifo_empty_tx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_3636_i_0_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_1_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_5), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(tx_dout_reg[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h599CC) )  un1_counter_cry_5_0 (.A(fifo_write_tx), 
        .B(fifo_read_tx), .C(\counter[5]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S_5), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_tx_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_2_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg({
        tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], tx_hold_reg[4], 
        tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], tx_hold_reg[0]})
        , .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_tx(fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(\counter[6]_net_1 ), 
        .FCI(un1_counter_cry_5), .S(un1_counter_s_6_S_5), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_304 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_304_FCO));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[5]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_2_fifo_256x8(
       tx_dout_reg,
       tx_hold_reg,
       fifo_write_tx,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_empty_tx,
       fifo_full_tx_i_0
    );
output [7:0] tx_dout_reg;
input  [7:0] tx_hold_reg;
input  fifo_write_tx;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_empty_tx;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_2_fifo_ctrl_128 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.tx_dout_reg({
        tx_dout_reg[7], tx_dout_reg[6], tx_dout_reg[5], tx_dout_reg[4], 
        tx_dout_reg[3], tx_dout_reg[2], tx_dout_reg[1], tx_dout_reg[0]})
        , .tx_hold_reg({tx_hold_reg[7], tx_hold_reg[6], tx_hold_reg[5], 
        tx_hold_reg[4], tx_hold_reg[3], tx_hold_reg[2], tx_hold_reg[1], 
        tx_hold_reg[0]}), .fifo_write_tx(fifo_write_tx), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    
endmodule


module mss_sb_CoreUARTapb_2_2_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       controlReg2,
       fifo_read_tx,
       fifo_read_tx_i_0,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       xmit_pulse_i_0,
       BT_RX_c,
       CoreUARTapb_2_2_TXRDY,
       fifo_full_tx_i_0,
       xmit_clock,
       baud_clock,
       fifo_empty_tx
    );
input  [7:0] tx_dout_reg;
input  [2:0] controlReg2;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  xmit_pulse_i_0;
output BT_RX_c;
output CoreUARTapb_2_2_TXRDY;
input  fifo_full_tx_i_0;
input  xmit_clock;
input  baud_clock;
input  fifo_empty_tx;

    wire \tx_byte[4]_net_1 , VCC_net_1, N_133_i_0, GND_net_1, 
        \tx_byte[5]_net_1 , \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_122_i_0, \xmit_bit_sel[2]_net_1 , 
        N_124_i_0, \xmit_bit_sel[3]_net_1 , N_126_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , \tx_byte[2]_net_1 , 
        \tx_byte[3]_net_1 , tx_parity_net_1, tx_parity_5, 
        un1_tx_parity_1_sqmuxa_0_1, tx_4_iv_i_0, N_144_i_0, 
        \xmit_state_ns_i_0[6] , \xmit_state[6]_net_1 , 
        \xmit_state_ns[6] , \xmit_state[0]_net_1 , 
        \xmit_state_ns[0]_net_1 , \xmit_state[1]_net_1 , 
        \xmit_state[2]_net_1 , \xmit_state_ns[2]_net_1 , 
        \xmit_state[3]_net_1 , N_112_i_0, \xmit_state[4]_net_1 , 
        \xmit_state_ns[4]_net_1 , \xmit_state[5]_net_1 , 
        \xmit_state_ns[5] , N_174, \xmit_state_ns_0_a2_2[5]_net_1 , 
        tx_2_u_i_m2_am_1_1, tx_2_u_i_m2_am_0, tx_2_u_i_m2_bm_1_1, 
        tx_2_u_i_m2_bm_0, N_487, N_377, N_413_1, N_408, 
        \xmit_state_ns_0_a2_3[5]_net_1 , N_172;
    
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(
        tx_2_u_i_m2_bm_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_bm_0));
    SLE tx_parity (.D(tx_parity_5), .CLK(GL0_INST), .EN(
        un1_tx_parity_1_sqmuxa_0_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(tx_parity_net_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(GL0_INST), .EN(VCC_net_1)
        , .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_2_TXRDY));
    CFG3 #( .INIT(8'hD8) )  \xmit_sel.tx_2_u_i_m2_ns  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(tx_2_u_i_m2_bm_0), .C(
        tx_2_u_i_m2_am_0), .Y(N_487));
    SLE \xmit_state[3]  (.D(N_112_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[3]_net_1 ));
    CFG3 #( .INIT(8'h82) )  \xmit_sel.tx_4_iv_0_a2  (.A(
        \xmit_state[4]_net_1 ), .B(controlReg2[2]), .C(tx_parity_net_1)
        , .Y(N_408));
    CFG4 #( .INIT(16'h0501) )  \xmit_sel.tx_4_iv_i  (.A(
        \xmit_state[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_408), 
        .D(N_487), .Y(tx_4_iv_i_0));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNI3UUF (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[4]_net_1 ));
    CFG4 #( .INIT(16'hFCAA) )  \xmit_state_ns_0[5]  (.A(
        \xmit_state[5]_net_1 ), .B(\xmit_state[4]_net_1 ), .C(
        \xmit_state_ns_0_a2_3[5]_net_1 ), .D(xmit_pulse_i_0), .Y(
        \xmit_state_ns[5] ));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3_0_a2[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_122_i_0));
    CFG2 #( .INIT(4'h7) )  \xmit_cnt.xmit_bit_sel_3_i_0_o2[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        N_377));
    VCC VCC (.Y(VCC_net_1));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[5]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_tx_parity_1_sqmuxa_0_a2_0_a2 (.A(
        \xmit_state[3]_net_1 ), .B(xmit_clock), .C(baud_clock), .D(
        controlReg2[1]), .Y(N_174));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_bm_1_1));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[5]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(
        xmit_pulse_i_0), .Y(\xmit_state_ns[2]_net_1 ));
    CFG4 #( .INIT(16'hAE0C) )  \xmit_state_ns[4]  (.A(N_172), .B(
        \xmit_state[4]_net_1 ), .C(xmit_pulse_i_0), .D(N_174), .Y(
        \xmit_state_ns[4]_net_1 ));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_126_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[3]_net_1 ));
    SLE \xmit_bit_sel[2]  (.D(N_124_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE tx (.D(tx_4_iv_i_0), .CLK(GL0_INST), .EN(N_144_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BT_RX_c));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[3]_net_1 ));
    CFG4 #( .INIT(16'h0804) )  \xmit_state_ns_i_a2_0_a2[3]  (.A(
        controlReg2[0]), .B(N_413_1), .C(\xmit_bit_sel[3]_net_1 ), .D(
        \xmit_bit_sel[0]_net_1 ), .Y(N_172));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[7]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_tx_parity_1_sqmuxa_0 (.A(N_174), .B(
        \xmit_state[5]_net_1 ), .Y(un1_tx_parity_1_sqmuxa_0_1));
    CFG4 #( .INIT(16'hF7C0) )  \xmit_state_RNO[3]  (.A(N_172), .B(
        xmit_pulse_i_0), .C(\xmit_state[2]_net_1 ), .D(
        \xmit_state[3]_net_1 ), .Y(N_112_i_0));
    CFG3 #( .INIT(8'h12) )  \xmit_par_calc.tx_parity_5  (.A(
        tx_parity_net_1), .B(\xmit_state[5]_net_1 ), .C(N_487), .Y(
        tx_parity_5));
    CFG2 #( .INIT(4'h8) )  \xmit_state_ns_0_a2_1[5]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[2]_net_1 ), .Y(
        N_413_1));
    CFG3 #( .INIT(8'h84) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(N_377), 
        .Y(N_124_i_0));
    CFG4 #( .INIT(16'h0400) )  \xmit_state_ns_0_a2_3[5]  (.A(
        controlReg2[1]), .B(\xmit_state_ns_0_a2_2[5]_net_1 ), .C(
        \xmit_bit_sel[3]_net_1 ), .D(\xmit_state[3]_net_1 ), .Y(
        \xmit_state_ns_0_a2_3[5]_net_1 ));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[6]_net_1 ));
    SLE \xmit_bit_sel[1]  (.D(N_122_i_0), .CLK(GL0_INST), .EN(
        xmit_pulse_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[1]_net_1 ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[1]_net_1 ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(GL0_INST), 
        .EN(xmit_pulse_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  fifo_read_en0_1_i_a3 (.A(fifo_empty_tx), .B(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[6] ));
    SLE fifo_read_en0 (.D(\xmit_state_ns_i_0[6] ), .CLK(GL0_INST), .EN(
        N_144_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_state_RNIH3M52[1]  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(
        xmit_pulse_i_0), .D(\xmit_state[6]_net_1 ), .Y(N_144_i_0));
    CFG2 #( .INIT(4'h8) )  \xmit_state_RNIKVA91[2]  (.A(xmit_pulse_i_0)
        , .B(\xmit_state[2]_net_1 ), .Y(N_133_i_0));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns[0]  (.A(fifo_empty_tx), 
        .B(xmit_pulse_i_0), .C(\xmit_state[5]_net_1 ), .D(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns[0]_net_1 ));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(GL0_INST), .EN(
        N_133_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \tx_byte[1]_net_1 ));
    SLE \xmit_state[4]  (.D(\xmit_state_ns[4]_net_1 ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\xmit_state[4]_net_1 ));
    CFG4 #( .INIT(16'hC600) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_bit_sel[3]_net_1 ), .C(
        N_377), .D(\xmit_state[3]_net_1 ), .Y(N_126_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_am_1_1));
    SLE \xmit_state[6]  (.D(\xmit_state_ns[6] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[6]_net_1 ));
    CFG2 #( .INIT(4'hB) )  fifo_read_en0_1_i_a3_i (.A(fifo_empty_tx), 
        .B(\xmit_state[0]_net_1 ), .Y(\xmit_state_ns_i_0[6] ));
    CFG4 #( .INIT(16'h8020) )  \xmit_state_ns_0_a2_2[5]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(controlReg2[0]), .Y(
        \xmit_state_ns_0_a2_2[5]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(
        tx_2_u_i_m2_am_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_am_0));
    
endmodule


module mss_sb_CoreUARTapb_2_2_Clock_gen_0s(
       controlReg1,
       controlReg2,
       xmit_clock,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       baud_clock,
       xmit_pulse_i_0
    );
input  [7:0] controlReg1;
input  [7:3] controlReg2;
output xmit_clock;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output baud_clock;
output xmit_pulse_i_0;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNI2H44_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIR89U2[8]  (.A(
        VCC_net_1), .B(controlReg2[3]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[8] ), .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] )
        , .Y(), .FCO(\baud_cntr_cry[8] ));
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[4] ));
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[1] ));
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[3] ));
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[3]_net_1 ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[9] ));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNI2H44  (.A(baud_cntr8_8)
        , .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(baud_cntr8_7), .FCI(
        VCC_net_1), .S(), .Y(baud_cntr8_1_RNI2H44_Y), .FCO(
        baud_cntr_cry_cy));
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNI2H44_Y), .CLK(
        GL0_INST), .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(baud_clock));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIUBTN[1]  (.A(
        VCC_net_1), .B(controlReg1[1]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[1] ), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] )
        , .Y(), .FCO(\baud_cntr_cry[1] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIQN3K3[10]  (.A(
        VCC_net_1), .B(controlReg2[5]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[10] ), .FCI(\baud_cntr_cry[9] ), .S(
        \baud_cntr_s[10] ), .Y(), .FCO(\baud_cntr_cry[10] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIFSP11[2]  (.A(
        VCC_net_1), .B(controlReg1[2]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[2] ), .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] )
        , .Y(), .FCO(\baud_cntr_cry[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI7JC92[6]  (.A(
        VCC_net_1), .B(controlReg1[6]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[6] ), .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] )
        , .Y(), .FCO(\baud_cntr_cry[6] ));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[7] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIM5993[9]  (.A(
        VCC_net_1), .B(controlReg2[4]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[9] ), .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] )
        , .Y(), .FCO(\baud_cntr_cry[9] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[5] ));
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[8] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI0CUU3[11]  (.A(
        VCC_net_1), .B(controlReg2[6]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[11] ), .FCI(\baud_cntr_cry[10] ), .S(
        \baud_cntr_s[11] ), .Y(), .FCO(\baud_cntr_cry[11] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIEQFV1[5]  (.A(
        VCC_net_1), .B(controlReg1[5]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[5] ), .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] )
        , .Y(), .FCO(\baud_cntr_cry[5] ));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[0] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI2FMB1[3]  (.A(
        VCC_net_1), .B(controlReg1[3]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[3] ), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] )
        , .Y(), .FCO(\baud_cntr_cry[3] ));
    CFG2 #( .INIT(4'h8) )  xmit_clock_RNI6E5R (.A(baud_clock), .B(
        xmit_clock), .Y(xmit_pulse_i_0));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNI2E9J2[7]  (.A(
        VCC_net_1), .B(controlReg1[7]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[7] ), .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] )
        , .Y(), .FCO(\baud_cntr_cry[7] ));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[10] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[6] ));
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(GL0_INST), .EN(
        baud_clock), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        xmit_clock));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h44700) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(controlReg2[7]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[12] ), .FCI(\baud_cntr_cry[11] ), .S(
        \baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[1]_net_1 ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIFT0E[0]  (.A(
        VCC_net_1), .B(controlReg1[0]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[0] ), .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), 
        .Y(), .FCO(\baud_cntr_cry[0] ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[2] ));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    ARI1 #( .INIT(20'h64700) )  \genblk1.baud_cntr_RNIN3JL1[4]  (.A(
        VCC_net_1), .B(controlReg1[4]), .C(baud_cntr8_1_RNI2H44_Y), .D(
        \baud_cntr[4] ), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] )
        , .Y(), .FCO(\baud_cntr_cry[4] ));
    
endmodule


module mss_sb_CoreUARTapb_2_2_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte_in,
       GL0_INST,
       MSS_HPMS_READY_int_RNI5CTC,
       fifo_write_rx_1
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte_in;
input  GL0_INST;
input  MSS_HPMS_READY_int_RNI5CTC;
input  fifo_write_rx_1;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(GL0_INST), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(MSS_HPMS_READY_int_RNI5CTC), 
        .A_DOUT_ARST_N(VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({
        rd_pointer[6], rd_pointer[5], rd_pointer[4], rd_pointer[3], 
        rd_pointer[2], rd_pointer[1], rd_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(
        VCC_net_1), .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(
        VCC_net_1), .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(
        VCC_net_1), .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(GL0_INST), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte_in[7], rx_byte_in[6], 
        rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], rx_byte_in[2], 
        rx_byte_in[1], rx_byte_in[0]}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_rx_1), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_2_fifo_ctrl_128_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_3652_i_0,
       N_3653_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_full_rx,
       fifo_empty_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_3652_i_0;
input  N_3653_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_full_rx;
output fifo_empty_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[1]_net_1 , VCC_net_1, 
        un1_counter_cry_1_0_S_6, GND_net_1, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_6, \counter[3]_net_1 , 
        un1_counter_cry_3_0_S_6, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_6, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_6, \counter[6]_net_1 , 
        un1_counter_s_6_S_6, \counter[0]_net_1 , un1_counter_cry_0_Y_5, 
        \data_out_0[0] , \data_out_0[1] , \data_out_0[2] , 
        \data_out_0[3] , \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \wr_pointer[1]_net_1 , 
        \wr_pointer_s[1] , \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_306_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_307_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_4_net_1, empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_307_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_2_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[2]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_1), 
        .S(un1_counter_cry_2_0_S_6), .Y(), .FCO(un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    SLE read_n_hold (.D(N_3652_i_0), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_4_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[4]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_3), 
        .S(un1_counter_cry_4_0_S_6), .Y(), .FCO(un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_306_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_306 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_306_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_6), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_3_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[3]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_2), 
        .S(un1_counter_cry_3_0_S_6), .Y(), .FCO(un1_counter_cry_3));
    ARI1 #( .INIT(20'h56699) )  un1_counter_cry_0 (.A(
        \counter[0]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(GND_net_1), .S(), .Y(
        un1_counter_cry_0_Y_5), .FCO(un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(\counter[0]_net_1 ), .B(
        empty_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_empty_rx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(GL0_INST), .EN(
        N_3653_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(GL0_INST), 
        .EN(fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_1_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[1]_net_1 ), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S_6), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNIIMDA (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(GL0_INST), .EN(
        read_n_hold_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout[1]));
    CFG4 #( .INIT(16'h8000) )  full (.A(\counter[0]_net_1 ), .B(
        full_4_net_1), .C(\counter[6]_net_1 ), .D(\counter[5]_net_1 ), 
        .Y(fifo_full_rx));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_307 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_307_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h566CC) )  un1_counter_cry_5_0 (.A(
        fifo_read_rx_0_sqmuxa), .B(fifo_write_rx_1), .C(
        \counter[5]_net_1 ), .D(GND_net_1), .FCI(un1_counter_cry_4), 
        .S(un1_counter_cry_5_0_S_6), .Y(), .FCO(un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(GL0_INST), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rd_pointer[4]_net_1 ));
    mss_sb_CoreUARTapb_2_2_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte_in({
        rx_byte_in[7], rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], 
        rx_byte_in[3], rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .GL0_INST(GL0_INST), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .fifo_write_rx_1(fifo_write_rx_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(
        \counter[6]_net_1 ), .FCI(un1_counter_cry_5), .S(
        un1_counter_s_6_S_6), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_5), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_4 (.A(\counter[4]_net_1 ), .B(
        \counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(full_4_net_1));
    
endmodule


module mss_sb_CoreUARTapb_2_2_fifo_256x8_0(
       rx_dout,
       rx_byte_in,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       N_3652_i_0,
       N_3653_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       fifo_full_rx,
       fifo_empty_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte_in;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  N_3652_i_0;
input  N_3653_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output fifo_full_rx;
output fifo_empty_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    mss_sb_CoreUARTapb_2_2_fifo_ctrl_128_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_byte_in({rx_byte_in[7], 
        rx_byte_in[6], rx_byte_in[5], rx_byte_in[4], rx_byte_in[3], 
        rx_byte_in[2], rx_byte_in[1], rx_byte_in[0]}), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_3652_i_0(N_3652_i_0), .N_3653_i_0(
        N_3653_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1), .fifo_full_rx(fifo_full_rx), 
        .fifo_empty_rx(fifo_empty_rx));
    
endmodule


module mss_sb_CoreUARTapb_2_2_COREUART_1s_1s_0s_15s_0s(
       CoreAPB3_0_APBmslave0_PWDATA,
       data_out,
       controlReg1,
       controlReg2,
       rx_dout_reg_5,
       rx_dout_reg_6,
       rx_dout_reg_7,
       rx_byte_7,
       rx_byte_6,
       rx_byte_5,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreUARTapb_2_2_OVERFLOW,
       CoreUARTapb_2_2_RXRDY,
       N_669,
       CoreAPB3_0_APBmslave4_PSELx,
       CoreUARTapb_2_2_PARITY_ERR,
       N_367,
       clear_overflow_0_a2_0_0,
       BT_RX_c,
       CoreUARTapb_2_2_TXRDY,
       BT_TX_c,
       CoreUARTapb_2_2_FRAMING_ERR
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [4:0] data_out;
input  [7:0] controlReg1;
input  [7:0] controlReg2;
output rx_dout_reg_5;
output rx_dout_reg_6;
output rx_dout_reg_7;
output rx_byte_7;
output rx_byte_6;
output rx_byte_5;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
output CoreUARTapb_2_2_OVERFLOW;
output CoreUARTapb_2_2_RXRDY;
input  N_669;
input  CoreAPB3_0_APBmslave4_PSELx;
output CoreUARTapb_2_2_PARITY_ERR;
input  N_367;
input  clear_overflow_0_a2_0_0;
output BT_RX_c;
output CoreUARTapb_2_2_TXRDY;
input  BT_TX_c;
output CoreUARTapb_2_2_FRAMING_ERR;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, 
        \rx_dout_reg[3]_net_1 , VCC_net_1, \rx_dout[3] , 
        rx_dout_reg4_i_0, GND_net_1, \rx_dout_reg[4]_net_1 , 
        \rx_dout[4] , \rx_dout[5] , \rx_dout[6] , \rx_dout[7] , 
        \tx_hold_reg[0]_net_1 , tx_hold_reg5, \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[4]_net_1 , \tx_hold_reg[5]_net_1 , 
        \tx_hold_reg[6]_net_1 , \tx_hold_reg[7]_net_1 , 
        \rx_dout_reg[0]_net_1 , \rx_dout[0] , \rx_dout_reg[1]_net_1 , 
        \rx_dout[1] , \rx_dout_reg[2]_net_1 , \rx_dout[2] , 
        \rx_state[0]_net_1 , \rx_state_ns[0] , \rx_state[1]_net_1 , 
        N_143_i, rx_dout_reg4, rx_dout_reg_empty_1_sqmuxa_i_0, 
        overflow_reg5_net_1, un1_clear_overflow_1, RXRDY5, 
        clear_parity_reg_net_1, clear_parity_reg0, clear_parity_en, 
        fifo_write_tx_net_1, tx_hold_reg5_i_0, fifo_empty_rx, 
        N_3652_i_0, fifo_full_rx, fifo_write, N_3653_i_0, \rx_byte[0] , 
        \rx_byte_in[0]_net_1 , \rx_byte[2] , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte[3] , \rx_byte_in[3]_net_1 , 
        \rx_byte[4] , \rx_byte_in[4]_net_1 , \rx_byte[1] , 
        \rx_byte_in[1]_net_1 , rx_idle, stop_strobe, 
        fifo_write_rx_1_net_1, fifo_read_rx_0_sqmuxa, xmit_clock, 
        baud_clock, xmit_pulse_i_0, \tx_dout_reg[0] , \tx_dout_reg[1] , 
        \tx_dout_reg[2] , \tx_dout_reg[3] , \tx_dout_reg[4] , 
        \tx_dout_reg[5] , \tx_dout_reg[6] , \tx_dout_reg[7] , 
        fifo_read_tx, fifo_read_tx_i_0, fifo_full_tx_i_0, 
        fifo_empty_tx;
    
    SLE \tx_hold_reg[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  overflow_reg5 (.A(fifo_full_rx), .B(
        fifo_write), .Y(overflow_reg5_net_1));
    CFG3 #( .INIT(8'h01) )  fifo_write_rx_1_i (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(N_3653_i_0));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[0]_net_1 ));
    CFG4 #( .INIT(16'hFFFB) )  fifo_read_rx_0_sqmuxa_0_a2_i (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(N_3652_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_143_i));
    CFG3 #( .INIT(8'hFE) )  fifo_write_rx_1 (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(fifo_full_rx), .C(fifo_write), 
        .Y(fifo_write_rx_1_net_1));
    mss_sb_CoreUARTapb_2_2_Rx_async_1s_0s_1s_2s make_RX (.rx_byte({
        rx_byte_7, rx_byte_6, rx_byte_5, \rx_byte[4] , \rx_byte[3] , 
        \rx_byte[2] , \rx_byte[1] , \rx_byte[0] }), .controlReg2({
        controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .clear_parity_reg(clear_parity_reg_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .BT_TX_c(BT_TX_c)
        , .CoreUARTapb_2_2_PARITY_ERR(CoreUARTapb_2_2_PARITY_ERR), 
        .stop_strobe(stop_strobe), .CoreUARTapb_2_2_FRAMING_ERR(
        CoreUARTapb_2_2_FRAMING_ERR), .clear_parity_en(clear_parity_en)
        , .fifo_write(fifo_write), .rx_idle(rx_idle));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[1]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\rx_byte[1] ), .Y(
        \rx_byte_in[1]_net_1 ));
    SLE \tx_hold_reg[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[3]_net_1 ));
    mss_sb_CoreUARTapb_2_2_fifo_256x8 \genblk2.tx_fifo  (.tx_dout_reg({
        \tx_dout_reg[7] , \tx_dout_reg[6] , \tx_dout_reg[5] , 
        \tx_dout_reg[4] , \tx_dout_reg[3] , \tx_dout_reg[2] , 
        \tx_dout_reg[1] , \tx_dout_reg[0] }), .tx_hold_reg({
        \tx_hold_reg[7]_net_1 , \tx_hold_reg[6]_net_1 , 
        \tx_hold_reg[5]_net_1 , \tx_hold_reg[4]_net_1 , 
        \tx_hold_reg[3]_net_1 , \tx_hold_reg[2]_net_1 , 
        \tx_hold_reg[1]_net_1 , \tx_hold_reg[0]_net_1 }), 
        .fifo_write_tx(fifo_write_tx_net_1), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_empty_tx(
        fifo_empty_tx), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[3]  (.A(\rx_byte[3] ), .B(
        CoreUARTapb_2_2_PARITY_ERR), .C(\rx_dout_reg[3]_net_1 ), .Y(
        data_out[3]));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE clear_framing_error_reg0 (.D(clear_parity_en), .CLK(GL0_INST), 
        .EN(VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(clear_parity_reg0));
    SLE \tx_hold_reg[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(GL0_INST), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(
        MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[5]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(rx_byte_5), .Y(
        \rx_byte_in[5]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  \genblk1.RXRDY5  (.A(rx_idle), .B(
        stop_strobe), .C(rx_dout_reg_empty_net_1), .Y(RXRDY5));
    CFG4 #( .INIT(16'h0004) )  fifo_read_rx_0_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(
        fifo_read_rx_0_sqmuxa));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[4]  (.A(\rx_byte[4] ), .B(
        CoreUARTapb_2_2_PARITY_ERR), .C(\rx_dout_reg[4]_net_1 ), .Y(
        data_out[4]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[2]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\rx_byte[2] ), .Y(
        \rx_byte_in[2]_net_1 ));
    mss_sb_CoreUARTapb_2_2_Tx_async_1s_0s_1s_2s_3s_4s_5s_6s make_TX (
        .tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .controlReg2({controlReg2[2], controlReg2[1], controlReg2[0]}), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .xmit_pulse_i_0(xmit_pulse_i_0), .BT_RX_c(BT_RX_c), 
        .CoreUARTapb_2_2_TXRDY(CoreUARTapb_2_2_TXRDY), 
        .fifo_full_tx_i_0(fifo_full_tx_i_0), .xmit_clock(xmit_clock), 
        .baud_clock(baud_clock), .fifo_empty_tx(fifo_empty_tx));
    SLE \tx_hold_reg[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[6]_net_1 ));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \reg_write.tx_hold_reg5_0_a2  (.A(N_669), 
        .B(CoreAPB3_0_APBmslave4_PSELx), .Y(tx_hold_reg5));
    mss_sb_CoreUARTapb_2_2_Clock_gen_0s make_CLOCK_GEN (.controlReg1({
        controlReg1[7], controlReg1[6], controlReg1[5], controlReg1[4], 
        controlReg1[3], controlReg1[2], controlReg1[1], controlReg1[0]})
        , .controlReg2({controlReg2[7], controlReg2[6], controlReg2[5], 
        controlReg2[4], controlReg2[3]}), .xmit_clock(xmit_clock), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .baud_clock(baud_clock), .xmit_pulse_i_0(
        xmit_pulse_i_0));
    SLE \rx_state[1]  (.D(N_143_i), .CLK(GL0_INST), .EN(VCC_net_1), 
        .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_7));
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[1]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  un1_clear_overflow (.A(N_367), .B(
        CoreAPB3_0_APBmslave4_PSELx), .C(overflow_reg5_net_1), .D(
        clear_overflow_0_a2_0_0), .Y(un1_clear_overflow_1));
    SLE clear_parity_reg (.D(clear_parity_reg0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        clear_parity_reg_net_1));
    CFG2 #( .INIT(4'h7) )  \reg_write.tx_hold_reg5_0_a2_i  (.A(N_669), 
        .B(CoreAPB3_0_APBmslave4_PSELx), .Y(tx_hold_reg5_i_0));
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_5));
    SLE overflow_reg (.D(overflow_reg5_net_1), .CLK(GL0_INST), .EN(
        un1_clear_overflow_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CoreUARTapb_2_2_OVERFLOW));
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[0]  (.A(\rx_byte[0] ), .B(
        CoreUARTapb_2_2_PARITY_ERR), .C(\rx_dout_reg[0]_net_1 ), .Y(
        data_out[0]));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[2]  (.A(\rx_byte[2] ), .B(
        CoreUARTapb_2_2_PARITY_ERR), .C(\rx_dout_reg[2]_net_1 ), .Y(
        data_out[2]));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_6));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \tx_hold_reg[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[7]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(GL0_INST), 
        .EN(RXRDY5), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreUARTapb_2_2_RXRDY));
    mss_sb_CoreUARTapb_2_2_fifo_256x8_0 \genblk3.rx_fifo  (.rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_byte_in({\rx_byte_in[7]_net_1 , \rx_byte_in[6]_net_1 , 
        \rx_byte_in[5]_net_1 , \rx_byte_in[4]_net_1 , 
        \rx_byte_in[3]_net_1 , \rx_byte_in[2]_net_1 , 
        \rx_byte_in[1]_net_1 , \rx_byte_in[0]_net_1 }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_3652_i_0(N_3652_i_0), .N_3653_i_0(
        N_3653_i_0), .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1_net_1), .fifo_full_rx(
        fifo_full_rx), .fifo_empty_rx(fifo_empty_rx));
    SLE \tx_hold_reg[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[3]_net_1 ));
    SLE fifo_write_tx (.D(tx_hold_reg5_i_0), .CLK(GL0_INST), .EN(
        VCC_net_1), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_write_tx_net_1));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[6]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(rx_byte_6), .Y(
        \rx_byte_in[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \DATA_OUT[1]  (.A(\rx_byte[1] ), .B(
        CoreUARTapb_2_2_PARITY_ERR), .C(\rx_dout_reg[1]_net_1 ), .Y(
        data_out[1]));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[7]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(rx_byte_7), .Y(
        \rx_byte_in[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[3]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\rx_byte[3] ), .Y(
        \rx_byte_in[3]_net_1 ));
    SLE \tx_hold_reg[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[1]_net_1 ));
    CFG4 #( .INIT(16'h8F0F) )  rx_dout_reg_empty_1_sqmuxa_i (.A(N_367), 
        .B(CoreAPB3_0_APBmslave4_PSELx), .C(rx_dout_reg4), .D(
        clear_overflow_0_a2_0_0), .Y(rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(GL0_INST), .EN(
        rx_dout_reg4_i_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\rx_dout_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[4]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\rx_byte[4] ), .Y(
        \rx_byte_in[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \rx_byte_in[0]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\rx_byte[0] ), .Y(
        \rx_byte_in[0]_net_1 ));
    SLE \tx_hold_reg[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(tx_hold_reg5), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\tx_hold_reg[4]_net_1 ));
    
endmodule


module 
        mss_sb_CoreUARTapb_2_2_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s(
        
       CoreAPB3_0_APBmslave0_PWDATA,
       CoreAPB3_0_APBmslave4_PRDATA,
       CoreAPB3_0_APBmslave0_PADDR,
       MSS_HPMS_READY_int_RNI5CTC,
       GL0_INST,
       CoreAPB3_0_APBmslave0_PWRITE,
       CoreAPB3_0_APBmslave0_PENABLE,
       N_437,
       CoreUARTapb_2_2_PARITY_ERR,
       N_99_1,
       psh_negedge_reg_1_sqmuxa_6_2,
       CoreAPB3_0_APBmslave4_PSELx,
       CoreUARTapb_2_2_TXRDY,
       CoreUARTapb_2_2_FRAMING_ERR,
       CoreUARTapb_2_2_OVERFLOW,
       CoreUARTapb_2_2_RXRDY,
       N_669,
       N_367,
       clear_overflow_0_a2_0_0,
       BT_RX_c,
       BT_TX_c
    );
input  [7:0] CoreAPB3_0_APBmslave0_PWDATA;
output [7:0] CoreAPB3_0_APBmslave4_PRDATA;
input  [4:2] CoreAPB3_0_APBmslave0_PADDR;
input  MSS_HPMS_READY_int_RNI5CTC;
input  GL0_INST;
input  CoreAPB3_0_APBmslave0_PWRITE;
input  CoreAPB3_0_APBmslave0_PENABLE;
output N_437;
output CoreUARTapb_2_2_PARITY_ERR;
input  N_99_1;
input  psh_negedge_reg_1_sqmuxa_6_2;
input  CoreAPB3_0_APBmslave4_PSELx;
output CoreUARTapb_2_2_TXRDY;
output CoreUARTapb_2_2_FRAMING_ERR;
output CoreUARTapb_2_2_OVERFLOW;
output CoreUARTapb_2_2_RXRDY;
input  N_669;
input  N_367;
input  clear_overflow_0_a2_0_0;
output BT_RX_c;
input  BT_TX_c;

    wire \controlReg1[4]_net_1 , VCC_net_1, controlReg14, GND_net_1, 
        \controlReg1[5]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[7]_net_1 , \NxtPrdata[5] , un1_NxtPrdata23_i_a2_0, 
        \NxtPrdata[6] , \NxtPrdata[7] , \controlReg2[0]_net_1 , 
        controlReg24, \controlReg2[1]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[7]_net_1 , \controlReg1[0]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[3]_net_1 , \NxtPrdata[0] , \NxtPrdata[1] , 
        \NxtPrdata[2] , \NxtPrdata[3] , \NxtPrdata[4] , 
        \NxtPrdata_5_bm_0[2] , \NxtPrdata_5_am_0[2] , 
        \NxtPrdata_5_bm_0[1] , \NxtPrdata_5_am_0[1] , 
        \NxtPrdata_5_bm[3]_net_1 , \NxtPrdata_5_am[3]_net_1 , 
        \NxtPrdata_5_bm[4]_net_1 , \NxtPrdata_5_am[4]_net_1 , 
        \NxtPrdata_5_bm[0]_net_1 , \NxtPrdata_5_am[0]_net_1 , 
        \NxtPrdata_5_bm[5]_net_1 , \NxtPrdata_5_am[5]_net_1 , 
        \NxtPrdata_5_bm[7]_net_1 , \NxtPrdata_5_am[7]_net_1 , 
        \NxtPrdata_5_bm[6]_net_1 , \NxtPrdata_5_am[6]_net_1 , 
        \rx_dout_reg[6] , \rx_byte[6] , \rx_dout_reg[7] , \rx_byte[7] , 
        \rx_dout_reg[5] , \rx_byte[5] , \data_out[0] , \data_out[4] , 
        \data_out[3] , \data_out[1] , \data_out[2] ;
    
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[4]  (.A(
        CoreUARTapb_2_2_FRAMING_ERR), .B(\data_out[4] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[4]_net_1 ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[5]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[5] ), 
        .D(\rx_byte[5] ), .Y(\NxtPrdata_5_am[5]_net_1 ));
    SLE \controlReg1[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[5]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[0]  (.A(
        CoreUARTapb_2_2_TXRDY), .B(\data_out[0] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[0]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[2]  (.A(
        \controlReg2[2]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[2]_net_1 ), .Y(\NxtPrdata_5_bm_0[2] ));
    SLE \controlReg1[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[7]_net_1 ));
    SLE \iPRDATA[1]  (.D(\NxtPrdata[1] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[1]));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[6]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[6] ), 
        .D(\rx_byte[6] ), .Y(\NxtPrdata_5_am[6]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[7]  (.A(
        \controlReg2[7]_net_1 ), .B(\controlReg1[7]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[7]_net_1 ));
    SLE \controlReg2[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[4]_net_1 ));
    SLE \iPRDATA[4]  (.D(\NxtPrdata[4] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[4]));
    CFG4 #( .INIT(16'h4000) )  \p_CtrlReg2Seq.controlReg24_0_a2_1  (.A(
        CoreAPB3_0_APBmslave0_PADDR[4]), .B(
        CoreAPB3_0_APBmslave0_PADDR[3]), .C(
        CoreAPB3_0_APBmslave0_PWRITE), .D(
        CoreAPB3_0_APBmslave0_PENABLE), .Y(N_437));
    VCC VCC (.Y(VCC_net_1));
    SLE \iPRDATA[3]  (.D(\NxtPrdata[3] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[3]));
    SLE \controlReg2[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[6]_net_1 ));
    SLE \controlReg1[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[4]  (.A(
        \controlReg2[4]_net_1 ), .B(\controlReg1[4]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[4]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[3]  (.A(
        CoreUARTapb_2_2_OVERFLOW), .B(\data_out[3] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[5]  (.A(
        \controlReg2[5]_net_1 ), .B(\controlReg1[5]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[5]_net_1 ));
    SLE \controlReg1[6]  (.D(CoreAPB3_0_APBmslave0_PWDATA[6]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[6]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[0]  (.A(
        \controlReg2[0]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[0]_net_1 ), .Y(\NxtPrdata_5_bm[0]_net_1 ));
    SLE \controlReg2[3]  (.D(CoreAPB3_0_APBmslave0_PWDATA[3]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[3]_net_1 ));
    SLE \controlReg1[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[2]_net_1 ));
    SLE \controlReg1[4]  (.D(CoreAPB3_0_APBmslave0_PWDATA[4]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[4]_net_1 ));
    SLE \iPRDATA[5]  (.D(\NxtPrdata[5] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[5]));
    SLE \iPRDATA[7]  (.D(\NxtPrdata[7] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[7]));
    SLE \controlReg2[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \p_CtrlReg2Seq.controlReg24_0_a2  (.A(
        CoreAPB3_0_APBmslave4_PSELx), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(controlReg24));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[6]  (.A(
        \controlReg2[6]_net_1 ), .B(\controlReg1[6]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[6]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[4]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[4]_net_1 ), 
        .C(\NxtPrdata_5_am[4]_net_1 ), .Y(\NxtPrdata[4] ));
    SLE \controlReg2[7]  (.D(CoreAPB3_0_APBmslave0_PWDATA[7]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[7]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[1]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[1] ), .C(
        \NxtPrdata_5_am_0[1] ), .Y(\NxtPrdata[1] ));
    SLE \iPRDATA[2]  (.D(\NxtPrdata[2] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[2]));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[0]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[0]_net_1 ), 
        .C(\NxtPrdata_5_am[0]_net_1 ), .Y(\NxtPrdata[0] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[3]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[3]_net_1 ), 
        .C(\NxtPrdata_5_am[3]_net_1 ), .Y(\NxtPrdata[3] ));
    SLE \controlReg2[5]  (.D(CoreAPB3_0_APBmslave0_PWDATA[5]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[5]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  \NxtPrdata_5_bm[3]  (.A(
        \controlReg2[3]_net_1 ), .B(\controlReg1[3]_net_1 ), .C(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_bm[3]_net_1 ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[1]  (.A(
        CoreUARTapb_2_2_RXRDY), .B(\data_out[1] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[1] ));
    SLE \controlReg2[2]  (.D(CoreAPB3_0_APBmslave0_PWDATA[2]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[2]_net_1 ));
    SLE \iPRDATA[6]  (.D(\NxtPrdata[6] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[6]));
    SLE \iPRDATA[0]  (.D(\NxtPrdata[0] ), .CLK(GL0_INST), .EN(
        un1_NxtPrdata23_i_a2_0), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CoreAPB3_0_APBmslave4_PRDATA[0]));
    mss_sb_CoreUARTapb_2_2_COREUART_1s_1s_0s_15s_0s uUART (
        .CoreAPB3_0_APBmslave0_PWDATA({CoreAPB3_0_APBmslave0_PWDATA[7], 
        CoreAPB3_0_APBmslave0_PWDATA[6], 
        CoreAPB3_0_APBmslave0_PWDATA[5], 
        CoreAPB3_0_APBmslave0_PWDATA[4], 
        CoreAPB3_0_APBmslave0_PWDATA[3], 
        CoreAPB3_0_APBmslave0_PWDATA[2], 
        CoreAPB3_0_APBmslave0_PWDATA[1], 
        CoreAPB3_0_APBmslave0_PWDATA[0]}), .data_out({\data_out[4] , 
        \data_out[3] , \data_out[2] , \data_out[1] , \data_out[0] }), 
        .controlReg1({\controlReg1[7]_net_1 , \controlReg1[6]_net_1 , 
        \controlReg1[5]_net_1 , \controlReg1[4]_net_1 , 
        \controlReg1[3]_net_1 , \controlReg1[2]_net_1 , 
        \controlReg1[1]_net_1 , \controlReg1[0]_net_1 }), .controlReg2({
        \controlReg2[7]_net_1 , \controlReg2[6]_net_1 , 
        \controlReg2[5]_net_1 , \controlReg2[4]_net_1 , 
        \controlReg2[3]_net_1 , \controlReg2[2]_net_1 , 
        \controlReg2[1]_net_1 , \controlReg2[0]_net_1 }), 
        .rx_dout_reg_5(\rx_dout_reg[5] ), .rx_dout_reg_6(
        \rx_dout_reg[6] ), .rx_dout_reg_7(\rx_dout_reg[7] ), 
        .rx_byte_7(\rx_byte[7] ), .rx_byte_6(\rx_byte[6] ), .rx_byte_5(
        \rx_byte[5] ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .CoreUARTapb_2_2_OVERFLOW(CoreUARTapb_2_2_OVERFLOW), 
        .CoreUARTapb_2_2_RXRDY(CoreUARTapb_2_2_RXRDY), .N_669(N_669), 
        .CoreAPB3_0_APBmslave4_PSELx(CoreAPB3_0_APBmslave4_PSELx), 
        .CoreUARTapb_2_2_PARITY_ERR(CoreUARTapb_2_2_PARITY_ERR), 
        .N_367(N_367), .clear_overflow_0_a2_0_0(
        clear_overflow_0_a2_0_0), .BT_RX_c(BT_RX_c), 
        .CoreUARTapb_2_2_TXRDY(CoreUARTapb_2_2_TXRDY), .BT_TX_c(
        BT_TX_c), .CoreUARTapb_2_2_FRAMING_ERR(
        CoreUARTapb_2_2_FRAMING_ERR));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[7]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[7]_net_1 ), 
        .C(\NxtPrdata_5_am[7]_net_1 ), .Y(\NxtPrdata[7] ));
    CFG4 #( .INIT(16'h0CA0) )  \NxtPrdata_5_am[2]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(\data_out[2] ), .C(
        CoreAPB3_0_APBmslave0_PADDR[4]), .D(
        CoreAPB3_0_APBmslave0_PADDR[2]), .Y(\NxtPrdata_5_am_0[2] ));
    SLE \controlReg2[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg24), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg2[0]_net_1 ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[2]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm_0[2] ), .C(
        \NxtPrdata_5_am_0[2] ), .Y(\NxtPrdata[2] ));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[6]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[6]_net_1 ), 
        .C(\NxtPrdata_5_am[6]_net_1 ), .Y(\NxtPrdata[6] ));
    CFG4 #( .INIT(16'hC840) )  \NxtPrdata_5_am[7]  (.A(
        CoreUARTapb_2_2_PARITY_ERR), .B(N_99_1), .C(\rx_dout_reg[7] ), 
        .D(\rx_byte[7] ), .Y(\NxtPrdata_5_am[7]_net_1 ));
    SLE \controlReg1[1]  (.D(CoreAPB3_0_APBmslave0_PWDATA[1]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[1]_net_1 ));
    CFG3 #( .INIT(8'h20) )  \p_CtrlReg1Seq.controlReg14_0_a2  (.A(
        CoreAPB3_0_APBmslave4_PSELx), .B(
        CoreAPB3_0_APBmslave0_PADDR[2]), .C(N_437), .Y(controlReg14));
    CFG3 #( .INIT(8'hB8) )  \NxtPrdata_5_bm[1]  (.A(
        \controlReg2[1]_net_1 ), .B(CoreAPB3_0_APBmslave0_PADDR[2]), 
        .C(\controlReg1[1]_net_1 ), .Y(\NxtPrdata_5_bm_0[1] ));
    CFG4 #( .INIT(16'h0100) )  un1_NxtPrdata23_i_a2 (.A(
        CoreAPB3_0_APBmslave0_PWRITE), .B(
        CoreAPB3_0_APBmslave0_PENABLE), .C(
        psh_negedge_reg_1_sqmuxa_6_2), .D(CoreAPB3_0_APBmslave4_PSELx), 
        .Y(un1_NxtPrdata23_i_a2_0));
    CFG3 #( .INIT(8'hD8) )  \NxtPrdata_5_ns[5]  (.A(
        CoreAPB3_0_APBmslave0_PADDR[3]), .B(\NxtPrdata_5_bm[5]_net_1 ), 
        .C(\NxtPrdata_5_am[5]_net_1 ), .Y(\NxtPrdata[5] ));
    SLE \controlReg1[0]  (.D(CoreAPB3_0_APBmslave0_PWDATA[0]), .CLK(
        GL0_INST), .EN(controlReg14), .ALn(MSS_HPMS_READY_int_RNI5CTC), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\controlReg1[0]_net_1 ));
    
endmodule


module mss_sb_CCC_0_FCCC(
       GL0_INST,
       LOCK_0,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output GL0_INST;
output LOCK_0;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST_inst_1 (.A(GL0_net), .Y(GL0_INST));
    CCC #( .INIT(210'h0000007FB8000045164000318C6318C1F18C61EC0404040400101)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        LOCK_0), .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(
        VCC_net_1), .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), 
        .NGMUX1_SEL(GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(
        GND_net_1), .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(
        VCC_net_1), .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(
        VCC_net_1), .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(
        VCC_net_1), .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(
        VCC_net_1), .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module mss_sb_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module mss_sb(
       PWM_c,
       COREI2C_0_0_SDA_IO,
       COREI2C_0_0_SCL_IO,
       DEVRST_N,
       mss_sb_0_TX,
       Echo_control_0_TX,
       GPS_RX_c,
       GPS_TX_c,
       BT_RX_c,
       BT_TX_c
    );
output [8:1] PWM_c;
inout  COREI2C_0_0_SDA_IO;
inout  COREI2C_0_0_SCL_IO;
input  DEVRST_N;
output mss_sb_0_TX;
input  Echo_control_0_TX;
output GPS_RX_c;
input  GPS_TX_c;
output BT_RX_c;
input  BT_TX_c;

    wire BIBUF_COREI2C_0_0_SDA_IO_Y, GND_net_1, 
        \COREI2C_0_0_SDAO_i[0] , BIBUF_COREI2C_0_0_SCL_IO_Y, 
        \COREI2C_0_0_SCLO_i[0] , SYSRESET_POR_net_1, 
        CoreUARTapb_2_2_intr_or_2_Y, CoreUARTapb_2_2_intr_or_1_Y, 
        CoreUARTapb_2_2_intr_or_0_Y, CoreUARTapb_2_2_RXRDY, 
        CoreUARTapb_2_2_TXRDY, CoreUARTapb_2_2_FRAMING_ERR, 
        CoreUARTapb_2_2_OVERFLOW, CoreUARTapb_2_2_PARITY_ERR, 
        CoreUARTapb_2_1_intr_or_2_Y, CoreUARTapb_2_1_intr_or_1_Y, 
        CoreUARTapb_2_1_intr_or_0_Y, CoreUARTapb_2_1_RXRDY, 
        CoreUARTapb_2_1_TXRDY, CoreUARTapb_2_1_FRAMING_ERR, 
        CoreUARTapb_2_1_OVERFLOW, CoreUARTapb_2_1_PARITY_ERR, 
        CoreUARTapb_2_0_intr_or_2_Y, CoreUARTapb_2_0_intr_or_1_Y, 
        CoreUARTapb_2_0_intr_or_0_Y, CoreUARTapb_2_0_RXRDY, 
        CoreUARTapb_2_0_TXRDY, CoreUARTapb_2_0_FRAMING_ERR, 
        CoreUARTapb_2_0_OVERFLOW, CoreUARTapb_2_0_PARITY_ERR, GL0_INST, 
        LOCK_0, FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] , \period_reg[5] , 
        \pwm_enable_reg[6] , \PRDATA_regif_0_0[5] , \sersta_m_0[1] , 
        \PRDATA_regif_9_i_0[4] , \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , \PRDATA_regif_9_i_1[4] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] , 
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \CoreAPB3_0_APBmslave4_PRDATA[2] , 
        \CoreAPB3_0_APBmslave4_PRDATA[3] , 
        \CoreAPB3_0_APBmslave4_PRDATA[4] , 
        \CoreAPB3_0_APBmslave4_PRDATA[5] , 
        \CoreAPB3_0_APBmslave4_PRDATA[6] , 
        \CoreAPB3_0_APBmslave4_PRDATA[7] , \serdat[4] , \serdat[0] , 
        \PRDATA_regif_12_0[1] , \PRDATAi[0][3] , \PRDATAi[0][1] , 
        \PRDATAi[0][7] , \PRDATAi[0][2] , \PRDATAi[0][5] , 
        \sersta_m[3] , \serdat_m[6] , \sercon_m[4] , \sercon_m[0] , 
        \sercon_m[6] , \CoreAPB3_0_APBmslave3_PRDATA[0] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PSELx, CoreAPB3_0_APBmslave4_PSELx, 
        CoreAPB3_0_APBmslave3_PSELx, CoreAPB3_0_APBmslave1_PSELx, 
        N_513, N_699, N_428, N_529, N_411, un12_PSELi, un9_PRDATA_2_0, 
        psh_enable_reg1_1_sqmuxa_0, N_629, N_432, N_685, N_680, N_684, 
        N_681, N_703, N_698, N_702, N_691, N_709, N_679, N_678, N_506, 
        N_711, N_140, N_710, un4_PRDATA, N_700, N_687, N_705, N_688, 
        N_706, N_690, N_708, N_689, N_707, N_686, N_704, 
        PRDATA_regif_sn_N_20_i_1, N_660, \COREI2C_0_0_INT[0] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , MSS_HPMS_READY_int_RNI5CTC, 
        N_528, CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, 
        \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[15] , 
        psh_negedge_reg_1_sqmuxa_6_2, N_425, N_423, 
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, N_99_1, N_367, N_437, 
        N_669, clear_overflow_0_a2_0_0, VCC_net_1;
    
    CoreAPB3_Z1_layer0 CoreAPB3_0 (
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] }), .period_reg({
        \period_reg[5] }), .pwm_enable_reg({\pwm_enable_reg[6] }), 
        .PRDATA_regif_0_0({\PRDATA_regif_0_0[5] }), .sersta_m_0({
        \sersta_m_0[1] }), .PRDATA_regif_9_i_0({
        \PRDATA_regif_9_i_0[4] }), .PRDATA_regif_9_i_1({
        \PRDATA_regif_9_i_1[4] }), .CoreAPB3_0_APBmslave4_PRDATA({
        \CoreAPB3_0_APBmslave4_PRDATA[7] , 
        \CoreAPB3_0_APBmslave4_PRDATA[6] , 
        \CoreAPB3_0_APBmslave4_PRDATA[5] , 
        \CoreAPB3_0_APBmslave4_PRDATA[4] , 
        \CoreAPB3_0_APBmslave4_PRDATA[3] , 
        \CoreAPB3_0_APBmslave4_PRDATA[2] , 
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] }), .PRDATA_regif_12_0({
        \PRDATA_regif_12_0[1] }), .sersta_m({\sersta_m[3] }), 
        .serdat_m({\serdat_m[6] }), .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PRDATA({
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR_3(
        \CoreAPB3_0_APBmslave0_PADDR[3] ), 
        .CoreAPB3_0_APBmslave0_PADDR_2(
        \CoreAPB3_0_APBmslave0_PADDR[2] ), 
        .CoreAPB3_0_APBmslave0_PADDR_0(
        \CoreAPB3_0_APBmslave0_PADDR[0] ), 
        .CoreAPB3_0_APBmslave0_PADDR_5(
        \CoreAPB3_0_APBmslave0_PADDR[5] ), .serdat_4(\serdat[4] ), 
        .serdat_0(\serdat[0] ), .\PRDATAi[0]_2 (\PRDATAi[0][3] ), 
        .\PRDATAi[0]_0 (\PRDATAi[0][1] ), .\PRDATAi[0]_6 (
        \PRDATAi[0][7] ), .\PRDATAi[0]_1 (\PRDATAi[0][2] ), 
        .\PRDATAi[0]_4 (\PRDATAi[0][5] ), .sercon_m_4(\sercon_m[4] ), 
        .sercon_m_0(\sercon_m[0] ), .sercon_m_6(\sercon_m[6] ), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave0_PSELx(CoreAPB3_0_APBmslave0_PSELx), 
        .CoreAPB3_0_APBmslave4_PSELx(CoreAPB3_0_APBmslave4_PSELx), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .N_513(N_513), .N_699(N_699), .N_428(N_428), .N_529(N_529), 
        .N_411(N_411), .un12_PSELi(un12_PSELi), .un9_PRDATA_2_0(
        un9_PRDATA_2_0), .psh_enable_reg1_1_sqmuxa_0(
        psh_enable_reg1_1_sqmuxa_0), .N_629(N_629), .N_432(N_432), 
        .N_685(N_685), .N_680(N_680), .N_684(N_684), .N_681(N_681), 
        .N_703(N_703), .N_698(N_698), .N_702(N_702), .N_691(N_691), 
        .N_709(N_709), .N_679(N_679), .N_678(N_678), .N_506(N_506), 
        .N_711(N_711), .N_140(N_140), .N_710(N_710), .un4_PRDATA(
        un4_PRDATA), .N_700(N_700), .N_687(N_687), .N_705(N_705), 
        .N_688(N_688), .N_706(N_706), .N_690(N_690), .N_708(N_708), 
        .N_689(N_689), .N_707(N_707), .N_686(N_686), .N_704(N_704), 
        .PRDATA_regif_sn_N_20_i_1(PRDATA_regif_sn_N_20_i_1), .N_660(
        N_660));
    BIBUF BIBUF_COREI2C_0_0_SDA_IO (.PAD(COREI2C_0_0_SDA_IO), .D(
        GND_net_1), .E(\COREI2C_0_0_SDAO_i[0] ), .Y(
        BIBUF_COREI2C_0_0_SDA_IO_Y));
    GND GND (.Y(GND_net_1));
    OR3 CoreUARTapb_2_1_intr_or_0 (.A(CoreUARTapb_2_1_FRAMING_ERR), .B(
        CoreUARTapb_2_1_OVERFLOW), .C(CoreUARTapb_2_1_PARITY_ERR), .Y(
        CoreUARTapb_2_1_intr_or_0_Y));
    OR3 CoreUARTapb_2_0_intr_or_1 (.A(CoreUARTapb_2_0_RXRDY), .B(
        CoreUARTapb_2_0_TXRDY), .C(GND_net_1), .Y(
        CoreUARTapb_2_0_intr_or_1_Y));
    COREI2C_Z2_layer0 COREI2C_0_0 (.COREI2C_0_0_SDAO_i({
        \COREI2C_0_0_SDAO_i[0] }), .COREI2C_0_0_SCLO_i({
        \COREI2C_0_0_SCLO_i[0] }), .COREI2C_0_0_INT({
        \COREI2C_0_0_INT[0] }), .CoreAPB3_0_APBmslave0_PADDR({
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] }), .sersta_m_0({
        \sersta_m_0[1] }), .sersta_m({\sersta_m[3] }), .serdat_m({
        \serdat_m[6] }), .CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .serdat_4(\serdat[4] ), 
        .serdat_0(\serdat[0] ), .sercon_m_6(\sercon_m[6] ), 
        .sercon_m_4(\sercon_m[4] ), .sercon_m_0(\sercon_m[0] ), 
        .\PRDATAi[0]_0 (\PRDATAi[0][1] ), .\PRDATAi[0]_1 (
        \PRDATAi[0][2] ), .\PRDATAi[0]_2 (\PRDATAi[0][3] ), 
        .\PRDATAi[0]_6 (\PRDATAi[0][7] ), .\PRDATAi[0]_4 (
        \PRDATAi[0][5] ), .un12_PSELi(un12_PSELi), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .un9_PRDATA_2_0(un9_PRDATA_2_0), 
        .BIBUF_COREI2C_0_0_SDA_IO_Y(BIBUF_COREI2C_0_0_SDA_IO_Y), 
        .BIBUF_COREI2C_0_0_SCL_IO_Y(BIBUF_COREI2C_0_0_SCL_IO_Y), 
        .N_528(N_528), .psh_enable_reg1_1_sqmuxa_0(
        psh_enable_reg1_1_sqmuxa_0), .un4_PRDATA(un4_PRDATA), 
        .CoreAPB3_0_APBmslave1_PSELx(CoreAPB3_0_APBmslave1_PSELx), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE));
    CoreResetP_Z6_layer0 CORERESETP_0 (.MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), 
        .SYSRESET_POR(SYSRESET_POR_net_1), 
        .mss_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), 
        .mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    OR3 CoreUARTapb_2_2_intr_or_1 (.A(CoreUARTapb_2_2_RXRDY), .B(
        CoreUARTapb_2_2_TXRDY), .C(GND_net_1), .Y(
        CoreUARTapb_2_2_intr_or_1_Y));
    OR3 CoreUARTapb_2_0_intr_or_2 (.A(CoreUARTapb_2_0_intr_or_1_Y), .B(
        CoreUARTapb_2_0_intr_or_0_Y), .C(GND_net_1), .Y(
        CoreUARTapb_2_0_intr_or_2_Y));
    OR3 CoreUARTapb_2_0_intr_or_0 (.A(CoreUARTapb_2_0_FRAMING_ERR), .B(
        CoreUARTapb_2_0_OVERFLOW), .C(CoreUARTapb_2_0_PARITY_ERR), .Y(
        CoreUARTapb_2_0_intr_or_0_Y));
    mss_sb_CoreUARTapb_2_0_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s 
        CoreUARTapb_2_0 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PRDATA({
        \CoreAPB3_0_APBmslave2_PRDATA[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_423(N_423), .N_99_1(N_99_1), .N_367(
        N_367), .CoreUARTapb_2_0_PARITY_ERR(CoreUARTapb_2_0_PARITY_ERR)
        , .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .psh_negedge_reg_1_sqmuxa_6_2(psh_negedge_reg_1_sqmuxa_6_2), 
        .N_432(N_432), .N_437(N_437), .CoreUARTapb_2_0_RXRDY(
        CoreUARTapb_2_0_RXRDY), .CoreUARTapb_2_0_TXRDY(
        CoreUARTapb_2_0_TXRDY), .CoreUARTapb_2_0_FRAMING_ERR(
        CoreUARTapb_2_0_FRAMING_ERR), .CoreUARTapb_2_0_OVERFLOW(
        CoreUARTapb_2_0_OVERFLOW), .N_669(N_669), 
        .clear_overflow_0_a2_0_0(clear_overflow_0_a2_0_0), 
        .mss_sb_0_TX(mss_sb_0_TX), .Echo_control_0_TX(
        Echo_control_0_TX));
    mss_sb_CoreUARTapb_2_1_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s 
        CoreUARTapb_2_1 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .N_425(N_425), .CoreUARTapb_2_1_OVERFLOW(
        CoreUARTapb_2_1_OVERFLOW), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .psh_negedge_reg_1_sqmuxa_6_2(
        psh_negedge_reg_1_sqmuxa_6_2), .CoreAPB3_0_APBmslave3_PSELx(
        CoreAPB3_0_APBmslave3_PSELx), .N_437(N_437), 
        .CoreUARTapb_2_1_PARITY_ERR(CoreUARTapb_2_1_PARITY_ERR), 
        .N_99_1(N_99_1), .N_367(N_367), .CoreUARTapb_2_1_FRAMING_ERR(
        CoreUARTapb_2_1_FRAMING_ERR), .CoreUARTapb_2_1_RXRDY(
        CoreUARTapb_2_1_RXRDY), .CoreUARTapb_2_1_TXRDY(
        CoreUARTapb_2_1_TXRDY), .N_669(N_669), 
        .clear_overflow_0_a2_0_0(clear_overflow_0_a2_0_0), .GPS_RX_c(
        GPS_RX_c), .GPS_TX_c(GPS_TX_c));
    OR3 CoreUARTapb_2_1_intr_or_2 (.A(CoreUARTapb_2_1_intr_or_1_Y), .B(
        CoreUARTapb_2_1_intr_or_0_Y), .C(GND_net_1), .Y(
        CoreUARTapb_2_1_intr_or_2_Y));
    corepwm_Z4_layer0 corepwm_0_0 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .PRDATA_regif_0_0({
        \PRDATA_regif_0_0[5] }), .CoreAPB3_0_APBmslave0_PADDR({
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), .PRDATA_regif_12_0({
        \PRDATA_regif_12_0[1] }), .PRDATA_regif_9_i_1({
        \PRDATA_regif_9_i_1[4] }), .PRDATA_regif_9_i_0({
        \PRDATA_regif_9_i_0[4] }), .PWM_c({PWM_c[8], PWM_c[7], 
        PWM_c[6], PWM_c[5], PWM_c[4], PWM_c[3], PWM_c[2], PWM_c[1]}), 
        .pwm_enable_reg_5(\pwm_enable_reg[6] ), .period_reg_5(
        \period_reg[5] ), .MSS_HPMS_READY_int_RNI5CTC(
        MSS_HPMS_READY_int_RNI5CTC), .GL0_INST(GL0_INST), .N_428(N_428)
        , .N_629(N_629), .N_678(N_678), .N_689(N_689), .N_686(N_686), 
        .N_679(N_679), .N_687(N_687), .N_688(N_688), .N_690(N_690), 
        .N_680(N_680), .N_685(N_685), .N_681(N_681), .N_684(N_684), 
        .N_691(N_691), .psh_enable_reg1_1_sqmuxa_0(
        psh_enable_reg1_1_sqmuxa_0), .N_528(N_528), 
        .psh_negedge_reg_1_sqmuxa_6_2(psh_negedge_reg_1_sqmuxa_6_2), 
        .N_529(N_529), .N_425(N_425), .N_423(N_423), .N_513(N_513), 
        .N_411(N_411), .N_660(N_660), .N_705(N_705), .N_706(N_706), 
        .N_708(N_708), .N_709(N_709), .N_711(N_711), .N_710(N_710), 
        .N_707(N_707), .N_704(N_704), .CoreAPB3_0_APBmslave0_PSELx(
        CoreAPB3_0_APBmslave0_PSELx), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .PRDATA_regif_sn_N_20_i_1(
        PRDATA_regif_sn_N_20_i_1), .N_506(N_506), .N_140(N_140), 
        .N_700(N_700), .N_702(N_702), .N_703(N_703), .N_699(N_699), 
        .N_698(N_698));
    mss_sb_MSS mss_sb_MSS_0 (.CoreAPB3_0_APBmslave0_PADDR({
        \CoreAPB3_0_APBmslave0_PADDR[8] , 
        \CoreAPB3_0_APBmslave0_PADDR[7] , 
        \CoreAPB3_0_APBmslave0_PADDR[6] , 
        \CoreAPB3_0_APBmslave0_PADDR[5] , 
        \CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] , 
        \CoreAPB3_0_APBmslave0_PADDR[1] , 
        \CoreAPB3_0_APBmslave0_PADDR[0] }), 
        .CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), .COREI2C_0_0_INT({
        \COREI2C_0_0_INT[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA({
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_3(
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[12] ), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_4(
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[13] ), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_5(
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[14] ), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR_6(
        \mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PADDR[15] ), 
        .mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        mss_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .CoreAPB3_0_APBmslave0_PENABLE(CoreAPB3_0_APBmslave0_PENABLE), 
        .mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx(
        mss_sb_MSS_TMP_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave0_PWRITE(CoreAPB3_0_APBmslave0_PWRITE), 
        .mss_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        mss_sb_MSS_TMP_0_MSS_RESET_N_M2F), 
        .CoreUARTapb_2_0_intr_or_2_Y(CoreUARTapb_2_0_intr_or_2_Y), 
        .CoreUARTapb_2_1_intr_or_2_Y(CoreUARTapb_2_1_intr_or_2_Y), 
        .CoreUARTapb_2_2_intr_or_2_Y(CoreUARTapb_2_2_intr_or_2_Y), 
        .LOCK_0(LOCK_0), .GL0_INST(GL0_INST));
    mss_sb_CoreUARTapb_2_2_CoreUARTapb_19s_1s_1s_1s_0s_0s_0s_0s_0s_0s 
        CoreUARTapb_2_2 (.CoreAPB3_0_APBmslave0_PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave4_PRDATA({
        \CoreAPB3_0_APBmslave4_PRDATA[7] , 
        \CoreAPB3_0_APBmslave4_PRDATA[6] , 
        \CoreAPB3_0_APBmslave4_PRDATA[5] , 
        \CoreAPB3_0_APBmslave4_PRDATA[4] , 
        \CoreAPB3_0_APBmslave4_PRDATA[3] , 
        \CoreAPB3_0_APBmslave4_PRDATA[2] , 
        \CoreAPB3_0_APBmslave4_PRDATA[1] , 
        \CoreAPB3_0_APBmslave4_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave0_PADDR({\CoreAPB3_0_APBmslave0_PADDR[4] , 
        \CoreAPB3_0_APBmslave0_PADDR[3] , 
        \CoreAPB3_0_APBmslave0_PADDR[2] }), 
        .MSS_HPMS_READY_int_RNI5CTC(MSS_HPMS_READY_int_RNI5CTC), 
        .GL0_INST(GL0_INST), .CoreAPB3_0_APBmslave0_PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .CoreAPB3_0_APBmslave0_PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .N_437(N_437), 
        .CoreUARTapb_2_2_PARITY_ERR(CoreUARTapb_2_2_PARITY_ERR), 
        .N_99_1(N_99_1), .psh_negedge_reg_1_sqmuxa_6_2(
        psh_negedge_reg_1_sqmuxa_6_2), .CoreAPB3_0_APBmslave4_PSELx(
        CoreAPB3_0_APBmslave4_PSELx), .CoreUARTapb_2_2_TXRDY(
        CoreUARTapb_2_2_TXRDY), .CoreUARTapb_2_2_FRAMING_ERR(
        CoreUARTapb_2_2_FRAMING_ERR), .CoreUARTapb_2_2_OVERFLOW(
        CoreUARTapb_2_2_OVERFLOW), .CoreUARTapb_2_2_RXRDY(
        CoreUARTapb_2_2_RXRDY), .N_669(N_669), .N_367(N_367), 
        .clear_overflow_0_a2_0_0(clear_overflow_0_a2_0_0), .BT_RX_c(
        BT_RX_c), .BT_TX_c(BT_TX_c));
    VCC VCC (.Y(VCC_net_1));
    OR3 CoreUARTapb_2_2_intr_or_0 (.A(CoreUARTapb_2_2_FRAMING_ERR), .B(
        CoreUARTapb_2_2_OVERFLOW), .C(CoreUARTapb_2_2_PARITY_ERR), .Y(
        CoreUARTapb_2_2_intr_or_0_Y));
    mss_sb_CCC_0_FCCC CCC_0 (.GL0_INST(GL0_INST), .LOCK_0(LOCK_0), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    BIBUF BIBUF_COREI2C_0_0_SCL_IO (.PAD(COREI2C_0_0_SCL_IO), .D(
        GND_net_1), .E(\COREI2C_0_0_SCLO_i[0] ), .Y(
        BIBUF_COREI2C_0_0_SCL_IO_Y));
    OR3 CoreUARTapb_2_2_intr_or_2 (.A(CoreUARTapb_2_2_intr_or_1_Y), .B(
        CoreUARTapb_2_2_intr_or_0_Y), .C(GND_net_1), .Y(
        CoreUARTapb_2_2_intr_or_2_Y));
    mss_sb_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    OR3 CoreUARTapb_2_1_intr_or_1 (.A(CoreUARTapb_2_1_RXRDY), .B(
        CoreUARTapb_2_1_TXRDY), .C(GND_net_1), .Y(
        CoreUARTapb_2_1_intr_or_1_Y));
    
endmodule


module pulse_meash(
       pulse_meash_0_tim,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       pulse_meash_0_new_ready,
       locator_control_0_en_timer,
       ECHO_c
    );
output [13:0] pulse_meash_0_tim;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
output pulse_meash_0_new_ready;
input  locator_control_0_en_timer;
input  ECHO_c;

    wire \i[9]_net_1 , \i_i[9] , \i[8]_net_1 , \i_i[8] , \i[7]_net_1 , 
        \i_i[7] , \i[6]_net_1 , \i_i[6] , \i[5]_net_1 , \i_i[5] , 
        \i[4]_net_1 , \i_i[4] , \i[15]_net_1 , \i_i[15] , 
        \i[14]_net_1 , \i_i[14] , \i[13]_net_1 , \i_i[13] , 
        \i[12]_net_1 , \i_i[12] , \i[11]_net_1 , \i_i[11] , 
        mult1_un152_sum_s_11_S, \mult1_un152_sum_i_0[13] , 
        mult1_un103_sum_s_11_S, \mult1_un103_sum_i_0[13] , 
        mult1_un110_sum_s_11_S, \mult1_un110_sum_i_0[13] , 
        mult1_un117_sum_s_11_S, \mult1_un117_sum_i_0[13] , 
        mult1_un124_sum_s_11_S, \mult1_un124_sum_i_0[13] , 
        mult1_un131_sum_s_11_S, \mult1_un131_sum_i_0[13] , 
        mult1_un138_sum_s_11_S, \mult1_un138_sum_i_0[13] , 
        mult1_un145_sum_s_11_S, \mult1_un145_sum_i_0[13] , 
        mult1_un68_sum_s_11_S, \mult1_un68_sum_i_0[13] , 
        mult1_un75_sum_s_11_S, \mult1_un75_sum_i_0[13] , 
        mult1_un82_sum_s_11_S, \mult1_un82_sum_i_0[13] , 
        mult1_un89_sum_s_11_S, \mult1_un89_sum_i_0[13] , 
        mult1_un96_sum_s_11_S, \mult1_un96_sum_i_0[13] , 
        mult1_un159_sum_s_11_S, \mult1_un159_sum_i_0[13] , VCC_net_1, 
        \state[1]_net_1 , GND_net_1, N_201_i_0, \state[0]_net_1 , 
        \state[4]_net_1 , N_183_i_0, \state[3]_net_1 , \state_ns[1] , 
        \state[2]_net_1 , N_5_i_0, N_187_i_0, \i[0]_net_1 , \i_s[0] , 
        \i[1]_net_1 , \i_s[1] , \i[2]_net_1 , \i_s[2] , \i[3]_net_1 , 
        \i_s[3] , \i_s[4] , \i_s[5] , \i_s[6] , \i_s[7] , \i_s[8] , 
        \i_s[9] , \i[10]_net_1 , \i_s[10] , \i_s[11] , \i_s[12] , 
        \i_s[13] , \i_s[14] , \i_s[15] , \i[16]_net_1 , \i_s[16] , 
        \i[17]_net_1 , \i_s[17] , \i[18]_net_1 , \i_s[18] , 
        \i[19]_net_1 , \i_s[19] , \i[20]_net_1 , \i_s[20] , CO2, 
        \i_s[21]_net_1 , \i_fast[19]_net_1 , \i_fast[20]_net_1 , 
        \i_fast[21]_net_1 , i_cry_cy, \i_cry[0]_net_1 , 
        \i_cry[1]_net_1 , \i_cry[2]_net_1 , \i_cry[3]_net_1 , 
        \i_cry[4]_net_1 , \i_cry[5]_net_1 , \i_cry[6]_net_1 , 
        \i_cry[7]_net_1 , \i_cry[8]_net_1 , \i_cry[9]_net_1 , 
        \i_cry[10]_net_1 , \i_cry[11]_net_1 , \i_cry[12]_net_1 , 
        \i_cry[13]_net_1 , \i_cry[14]_net_1 , \i_cry[15]_net_1 , 
        \i_cry[16]_net_1 , \i_cry[17]_net_1 , \i_cry[18]_net_1 , 
        \i_cry[19]_net_1 , \i_cry[20]_net_1 , mult1_un159_sum_cry_0, 
        mult1_un159_sum_cry_1, mult1_un152_sum_cry_0_Y, 
        mult1_un159_sum_cry_2, mult1_un152_sum_cry_1_S, 
        mult1_un159_sum_cry_3, mult1_un152_sum_cry_2_S, 
        mult1_un159_sum_cry_4, mult1_un152_sum_cry_3_S, 
        mult1_un159_sum_cry_5, mult1_un152_sum_cry_4_S, 
        mult1_un159_sum_cry_6, mult1_un152_sum_cry_5_S, 
        mult1_un159_sum_cry_7, mult1_un152_sum_cry_6_S, 
        mult1_un159_sum_cry_8, mult1_un152_sum_cry_7_S, 
        mult1_un159_sum_cry_9, mult1_un152_sum_cry_8_S, 
        mult1_un152_sum_cry_10_S, mult1_un159_sum_cry_10, 
        mult1_un152_sum_cry_9_S, mult1_un110_sum_cry_0, 
        mult1_un110_sum_cry_1, mult1_un110_sum_cry_1_S, 
        mult1_un103_sum_cry_0_Y, mult1_un110_sum_cry_2, 
        mult1_un110_sum_cry_2_S, mult1_un103_sum_cry_1_S, 
        mult1_un110_sum_cry_3, mult1_un110_sum_cry_3_S, 
        mult1_un103_sum_cry_2_S, mult1_un110_sum_cry_4, 
        mult1_un110_sum_cry_4_S, mult1_un103_sum_cry_3_S, 
        mult1_un110_sum_cry_5, mult1_un110_sum_cry_5_S, 
        mult1_un103_sum_cry_4_S, mult1_un110_sum_cry_6, 
        mult1_un110_sum_cry_6_S, mult1_un103_sum_cry_5_S, 
        mult1_un110_sum_cry_7, mult1_un110_sum_cry_7_S, 
        mult1_un103_sum_cry_6_S, mult1_un110_sum_cry_8, 
        mult1_un110_sum_cry_8_S, mult1_un103_sum_cry_7_S, 
        mult1_un110_sum_cry_9, mult1_un110_sum_cry_9_S, 
        mult1_un103_sum_cry_8_S, mult1_un103_sum_cry_10_S, 
        mult1_un110_sum_cry_10, mult1_un110_sum_cry_10_S, 
        mult1_un103_sum_cry_9_S, mult1_un117_sum_cry_0, 
        mult1_un117_sum_cry_1, mult1_un117_sum_cry_1_S, 
        mult1_un117_sum_cry_2, mult1_un117_sum_cry_2_S, 
        mult1_un117_sum_cry_3, mult1_un117_sum_cry_3_S, 
        mult1_un117_sum_cry_4, mult1_un117_sum_cry_4_S, 
        mult1_un117_sum_cry_5, mult1_un117_sum_cry_5_S, 
        mult1_un117_sum_cry_6, mult1_un117_sum_cry_6_S, 
        mult1_un117_sum_cry_7, mult1_un117_sum_cry_7_S, 
        mult1_un117_sum_cry_8, mult1_un117_sum_cry_8_S, 
        mult1_un117_sum_cry_9, mult1_un117_sum_cry_9_S, 
        mult1_un117_sum_cry_10, mult1_un117_sum_cry_10_S, 
        mult1_un124_sum_cry_0, mult1_un124_sum_cry_1, 
        mult1_un124_sum_cry_1_S, mult1_un124_sum_cry_2, 
        mult1_un124_sum_cry_2_S, mult1_un124_sum_cry_3, 
        mult1_un124_sum_cry_3_S, mult1_un124_sum_cry_4, 
        mult1_un124_sum_cry_4_S, mult1_un124_sum_cry_5, 
        mult1_un124_sum_cry_5_S, mult1_un124_sum_cry_6, 
        mult1_un124_sum_cry_6_S, mult1_un124_sum_cry_7, 
        mult1_un124_sum_cry_7_S, mult1_un124_sum_cry_8, 
        mult1_un124_sum_cry_8_S, mult1_un124_sum_cry_9, 
        mult1_un124_sum_cry_9_S, mult1_un124_sum_cry_10, 
        mult1_un124_sum_cry_10_S, mult1_un131_sum_cry_0, 
        mult1_un131_sum_cry_1, mult1_un131_sum_cry_1_S, 
        mult1_un131_sum_cry_2, mult1_un131_sum_cry_2_S, 
        mult1_un131_sum_cry_3, mult1_un131_sum_cry_3_S, 
        mult1_un131_sum_cry_4, mult1_un131_sum_cry_4_S, 
        mult1_un131_sum_cry_5, mult1_un131_sum_cry_5_S, 
        mult1_un131_sum_cry_6, mult1_un131_sum_cry_6_S, 
        mult1_un131_sum_cry_7, mult1_un131_sum_cry_7_S, 
        mult1_un131_sum_cry_8, mult1_un131_sum_cry_8_S, 
        mult1_un131_sum_cry_9, mult1_un131_sum_cry_9_S, 
        mult1_un131_sum_cry_10, mult1_un131_sum_cry_10_S, 
        mult1_un138_sum_cry_0, mult1_un138_sum_cry_1, 
        mult1_un138_sum_cry_1_S, mult1_un138_sum_cry_2, 
        mult1_un138_sum_cry_2_S, mult1_un138_sum_cry_3, 
        mult1_un138_sum_cry_3_S, mult1_un138_sum_cry_4, 
        mult1_un138_sum_cry_4_S, mult1_un138_sum_cry_5, 
        mult1_un138_sum_cry_5_S, mult1_un138_sum_cry_6, 
        mult1_un138_sum_cry_6_S, mult1_un138_sum_cry_7, 
        mult1_un138_sum_cry_7_S, mult1_un138_sum_cry_8, 
        mult1_un138_sum_cry_8_S, mult1_un138_sum_cry_9, 
        mult1_un138_sum_cry_9_S, mult1_un138_sum_cry_10, 
        mult1_un138_sum_cry_10_S, mult1_un145_sum_cry_0, 
        mult1_un145_sum_cry_1, mult1_un145_sum_cry_1_S, 
        mult1_un145_sum_cry_2, mult1_un145_sum_cry_2_S, 
        mult1_un145_sum_cry_3, mult1_un145_sum_cry_3_S, 
        mult1_un145_sum_cry_4, mult1_un145_sum_cry_4_S, 
        mult1_un145_sum_cry_5, mult1_un145_sum_cry_5_S, 
        mult1_un145_sum_cry_6, mult1_un145_sum_cry_6_S, 
        mult1_un145_sum_cry_7, mult1_un145_sum_cry_7_S, 
        mult1_un145_sum_cry_8, mult1_un145_sum_cry_8_S, 
        mult1_un145_sum_cry_9, mult1_un145_sum_cry_9_S, 
        mult1_un145_sum_cry_10, mult1_un145_sum_cry_10_S, 
        mult1_un152_sum_cry_0, mult1_un152_sum_cry_1, 
        mult1_un152_sum_cry_2, mult1_un152_sum_cry_3, 
        mult1_un152_sum_cry_4, mult1_un152_sum_cry_5, 
        mult1_un152_sum_cry_6, mult1_un152_sum_cry_7, 
        mult1_un152_sum_cry_8, mult1_un152_sum_cry_9, 
        mult1_un152_sum_cry_10, mult1_un54_sum_cry_0, 
        mult1_un54_sum_cry_1, mult1_un54_sum_cry_1_S, 
        mult1_un47_sum_cry_0_Y, mult1_un54_sum_cry_2, 
        mult1_un61_sum_axb_3, mult1_un47_sum_cry_1_S, 
        mult1_un54_sum_cry_3, mult1_un54_sum_cry_3_S, 
        mult1_un54_sum_axb_3, mult1_un54_sum_cry_4, 
        mult1_un61_sum_axb_5, mult1_un47_sum_cry_3_S, 
        mult1_un54_sum_cry_5, mult1_un54_sum_cry_5_S, 
        mult1_un54_sum_axb_5, mult1_un54_sum_cry_6, 
        mult1_un54_sum_cry_6_S, mult1_un47_sum_s_5_sf, 
        mult1_un47_sum_cry_4, mult1_un54_sum_s_8_S, 
        mult1_un54_sum_cry_7, mult1_un61_sum_axb_8, 
        mult1_un61_sum_cry_0, mult1_un61_sum_cry_1, 
        mult1_un61_sum_cry_1_S, mult1_un61_sum_cry_2, 
        mult1_un68_sum_axb_3, mult1_un61_sum_cry_3, 
        mult1_un61_sum_cry_3_S, mult1_un61_sum_cry_4, 
        mult1_un68_sum_axb_5, mult1_un61_sum_cry_5, 
        mult1_un61_sum_cry_5_S, mult1_un61_sum_cry_6, 
        mult1_un61_sum_cry_6_S, mult1_un61_sum_cry_7, 
        mult1_un68_sum_axb_8, mult1_un61_sum_cry_8, 
        mult1_un61_sum_cry_8_S, mult1_un68_sum_axb_11, 
        mult1_un61_sum_cry_9, mult1_un68_sum_axb_10, 
        mult1_un68_sum_cry_0, mult1_un68_sum_cry_1, 
        mult1_un68_sum_cry_1_S, mult1_un68_sum_cry_2, 
        mult1_un68_sum_cry_2_S, mult1_un68_sum_cry_3, 
        mult1_un68_sum_cry_3_S, mult1_un68_sum_cry_4, 
        mult1_un68_sum_cry_4_S, mult1_un68_sum_cry_5, 
        mult1_un68_sum_cry_5_S, mult1_un68_sum_cry_6, 
        mult1_un68_sum_cry_6_S, mult1_un68_sum_cry_7, 
        mult1_un68_sum_cry_7_S, mult1_un68_sum_cry_8, 
        mult1_un68_sum_cry_8_S, mult1_un68_sum_cry_9, 
        mult1_un68_sum_cry_9_S, mult1_un68_sum_cry_10, 
        mult1_un68_sum_cry_10_S, mult1_un75_sum_cry_0, 
        mult1_un75_sum_cry_1, mult1_un75_sum_cry_1_S, 
        mult1_un75_sum_cry_2, mult1_un75_sum_cry_2_S, 
        mult1_un75_sum_cry_3, mult1_un75_sum_cry_3_S, 
        mult1_un75_sum_cry_4, mult1_un75_sum_cry_4_S, 
        mult1_un75_sum_cry_5, mult1_un75_sum_cry_5_S, 
        mult1_un75_sum_cry_6, mult1_un75_sum_cry_6_S, 
        mult1_un75_sum_cry_7, mult1_un75_sum_cry_7_S, 
        mult1_un75_sum_cry_8, mult1_un75_sum_cry_8_S, 
        mult1_un75_sum_cry_9, mult1_un75_sum_cry_9_S, 
        mult1_un75_sum_cry_10, mult1_un75_sum_cry_10_S, 
        mult1_un82_sum_cry_0, mult1_un82_sum_cry_1, 
        mult1_un82_sum_cry_1_S, mult1_un82_sum_cry_2, 
        mult1_un82_sum_cry_2_S, mult1_un82_sum_cry_3, 
        mult1_un82_sum_cry_3_S, mult1_un82_sum_cry_4, 
        mult1_un82_sum_cry_4_S, mult1_un82_sum_cry_5, 
        mult1_un82_sum_cry_5_S, mult1_un82_sum_cry_6, 
        mult1_un82_sum_cry_6_S, mult1_un82_sum_cry_7, 
        mult1_un82_sum_cry_7_S, mult1_un82_sum_cry_8, 
        mult1_un82_sum_cry_8_S, mult1_un82_sum_cry_9, 
        mult1_un82_sum_cry_9_S, mult1_un82_sum_cry_10, 
        mult1_un82_sum_cry_10_S, mult1_un89_sum_cry_0, 
        mult1_un89_sum_cry_1, mult1_un89_sum_cry_1_S, 
        mult1_un89_sum_cry_2, mult1_un89_sum_cry_2_S, 
        mult1_un89_sum_cry_3, mult1_un89_sum_cry_3_S, 
        mult1_un89_sum_cry_4, mult1_un89_sum_cry_4_S, 
        mult1_un89_sum_cry_5, mult1_un89_sum_cry_5_S, 
        mult1_un89_sum_cry_6, mult1_un89_sum_cry_6_S, 
        mult1_un89_sum_cry_7, mult1_un89_sum_cry_7_S, 
        mult1_un89_sum_cry_8, mult1_un89_sum_cry_8_S, 
        mult1_un89_sum_cry_9, mult1_un89_sum_cry_9_S, 
        mult1_un89_sum_cry_10, mult1_un89_sum_cry_10_S, 
        mult1_un96_sum_cry_0, mult1_un96_sum_cry_1, 
        mult1_un96_sum_cry_1_S, mult1_un96_sum_cry_2, 
        mult1_un96_sum_cry_2_S, mult1_un96_sum_cry_3, 
        mult1_un96_sum_cry_3_S, mult1_un96_sum_cry_4, 
        mult1_un96_sum_cry_4_S, mult1_un96_sum_cry_5, 
        mult1_un96_sum_cry_5_S, mult1_un96_sum_cry_6, 
        mult1_un96_sum_cry_6_S, mult1_un96_sum_cry_7, 
        mult1_un96_sum_cry_7_S, mult1_un96_sum_cry_8, 
        mult1_un96_sum_cry_8_S, mult1_un96_sum_cry_9, 
        mult1_un96_sum_cry_9_S, mult1_un96_sum_cry_10, 
        mult1_un96_sum_cry_10_S, mult1_un103_sum_cry_0, 
        mult1_un103_sum_cry_1, mult1_un103_sum_cry_2, 
        mult1_un103_sum_cry_3, mult1_un103_sum_cry_4, 
        mult1_un103_sum_cry_5, mult1_un103_sum_cry_6, 
        mult1_un103_sum_cry_7, mult1_un103_sum_cry_8, 
        mult1_un103_sum_cry_9, mult1_un103_sum_cry_10, 
        mult1_un47_sum_cry_0, mult1_un47_sum_cry_1, 
        mult1_un47_sum_cry_2, mult1_un47_sum_cry_3, 
        \state_ns_i_0_0[0]_net_1 , un20_clklto16_1_net_1, un20_clklt9, 
        un20_clklt12, un20_clklt16, un20_clklt20, 
        \state_ns_o2[2]_net_1 ;
    
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_1  (.A(\i_i[14] ), 
        .B(mult1_un75_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un82_sum_cry_0), .S(mult1_un82_sum_cry_1_S), .Y(), .FCO(
        mult1_un82_sum_cry_1));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_9  (.A(
        mult1_un89_sum_cry_8_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_8), .S(
        mult1_un96_sum_cry_9_S), .Y(), .FCO(mult1_un96_sum_cry_9));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_5  (.A(
        mult1_un124_sum_cry_4_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_4), .S(
        mult1_un131_sum_cry_5_S), .Y(), .FCO(mult1_un131_sum_cry_5));
    SLE \state[0]  (.D(\state[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \i_RNI4BK2[4]  (.A(\i[4]_net_1 ), .Y(
        \i_i[4] ));
    ARI1 #( .INIT(20'h45500) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_cry_1  (.A(VCC_net_1), 
        .B(\i_fast[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un47_sum_cry_0), .S(mult1_un47_sum_cry_1_S), .Y(), .FCO(
        mult1_un47_sum_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_1  (.A(\i_i[8] ), 
        .B(mult1_un117_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un124_sum_cry_0), .S(mult1_un124_sum_cry_1_S), .Y(), 
        .FCO(mult1_un124_sum_cry_1));
    SLE \i[7]  (.D(\i_s[7] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_i_0[13]  (.A(
        mult1_un89_sum_s_11_S), .Y(\mult1_un89_sum_i_0[13] ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_i_0[13]  (.A(
        mult1_un110_sum_s_11_S), .Y(\mult1_un110_sum_i_0[13] ));
    SLE \i[16]  (.D(\i_s[16] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[16]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_3  (.A(
        mult1_un145_sum_cry_2_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_2), .S(
        mult1_un152_sum_cry_3_S), .Y(), .FCO(mult1_un152_sum_cry_3));
    ARI1 #( .INIT(20'h42200) )  \i_s[21]  (.A(VCC_net_1), .B(CO2), .C(
        \state[3]_net_1 ), .D(GND_net_1), .FCI(\i_cry[20]_net_1 ), .S(
        \i_s[21]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_5  (.A(
        mult1_un68_sum_cry_4_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_4), .S(
        mult1_un75_sum_cry_5_S), .Y(), .FCO(mult1_un75_sum_cry_5));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un159_sum_cry_0));
    SLE \tim[4]  (.D(\mult1_un131_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[4]));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_i_0[13]  (.A(
        mult1_un124_sum_s_11_S), .Y(\mult1_un124_sum_i_0[13] ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[14]  (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[13]_net_1 ), .S(\i_s[14] ), .Y(), .FCO(
        \i_cry[14]_net_1 ));
    ARI1 #( .INIT(20'h6E000) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_cry_4  (.A(VCC_net_1), 
        .B(\i_fast[19]_net_1 ), .C(\i_fast[20]_net_1 ), .D(
        \i_fast[21]_net_1 ), .FCI(mult1_un47_sum_cry_3), .S(
        mult1_un54_sum_axb_5), .Y(), .FCO(mult1_un47_sum_cry_4));
    SLE \i[21]  (.D(\i_s[21]_net_1 ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(CO2));
    ARI1 #( .INIT(20'h42200) )  \i_cry[20]  (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[19]_net_1 ), .S(\i_s[20] ), .Y(), .FCO(
        \i_cry[20]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_3  (.A(
        mult1_un82_sum_cry_2_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_2), .S(
        mult1_un89_sum_cry_3_S), .Y(), .FCO(mult1_un89_sum_cry_3));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un89_sum_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_8  (.A(
        mult1_un131_sum_cry_7_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_7), .S(
        mult1_un138_sum_cry_8_S), .Y(), .FCO(mult1_un138_sum_cry_8));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_8  (.A(VCC_net_1), 
        .B(mult1_un61_sum_axb_8), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_7), .S(mult1_un61_sum_cry_8_S), .Y(), .FCO(
        mult1_un61_sum_cry_8));
    SLE \i[0]  (.D(\i_s[0] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_7  (.A(
        mult1_un89_sum_cry_6_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_6), .S(
        mult1_un96_sum_cry_7_S), .Y(), .FCO(mult1_un96_sum_cry_7));
    SLE \i[11]  (.D(\i_s[11] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(mult1_un152_sum_cry_0_Y), .FCO(
        mult1_un152_sum_cry_0));
    CFG2 #( .INIT(4'hE) )  \state_ns_i_0_0[0]  (.A(\state[3]_net_1 ), 
        .B(\state[2]_net_1 ), .Y(\state_ns_i_0_0[0]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_3  (.A(
        mult1_un89_sum_cry_2_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_2), .S(
        mult1_un96_sum_cry_3_S), .Y(), .FCO(mult1_un96_sum_cry_3));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_2  (.A(
        mult1_un82_sum_cry_1_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_1), .S(
        mult1_un89_sum_cry_2_S), .Y(), .FCO(mult1_un89_sum_cry_2));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_4  (.A(
        mult1_un138_sum_cry_3_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_3), .S(
        mult1_un145_sum_cry_4_S), .Y(), .FCO(mult1_un145_sum_cry_4));
    ARI1 #( .INIT(20'h55555) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_1  (.A(VCC_net_1), 
        .B(\i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_0), .S(mult1_un61_sum_cry_1_S), .Y(), .FCO(
        mult1_un61_sum_cry_1));
    CFG3 #( .INIT(8'h4F) )  \state_ns_o2_3[2]  (.A(\i[9]_net_1 ), .B(
        un20_clklt9), .C(\i[10]_net_1 ), .Y(un20_clklt12));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_10  (.A(VCC_net_1)
        , .B(mult1_un68_sum_axb_10), .C(GND_net_1), .D(GND_net_1), 
        .FCI(mult1_un68_sum_cry_9), .S(mult1_un68_sum_cry_10_S), .Y(), 
        .FCO(mult1_un68_sum_cry_10));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_10  (.A(
        mult1_un138_sum_cry_9_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_9), .S(
        mult1_un145_sum_cry_10_S), .Y(), .FCO(mult1_un145_sum_cry_10));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_4  (.A(
        mult1_un124_sum_cry_3_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_3), .S(
        mult1_un131_sum_cry_4_S), .Y(), .FCO(mult1_un131_sum_cry_4));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_2  (.A(VCC_net_1), 
        .B(mult1_un61_sum_cry_1_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_1), .S(mult1_un68_sum_cry_2_S), .Y(), .FCO(
        mult1_un68_sum_cry_2));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_4  (.A(
        mult1_un96_sum_cry_3_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_3), .S(
        mult1_un103_sum_cry_4_S), .Y(), .FCO(mult1_un103_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_9  (.A(
        mult1_un117_sum_cry_8_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_8), .S(
        mult1_un124_sum_cry_9_S), .Y(), .FCO(mult1_un124_sum_cry_9));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_4  (.A(
        mult1_un89_sum_cry_3_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_3), .S(
        mult1_un96_sum_cry_4_S), .Y(), .FCO(mult1_un96_sum_cry_4));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_1  (.A(\i_i[9] ), 
        .B(mult1_un110_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un117_sum_cry_0), .S(mult1_un117_sum_cry_1_S), .Y(), 
        .FCO(mult1_un117_sum_cry_1));
    ARI1 #( .INIT(20'h66600) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_cry_2  (.A(VCC_net_1), 
        .B(\i_fast[19]_net_1 ), .C(\i_fast[20]_net_1 ), .D(GND_net_1), 
        .FCI(mult1_un47_sum_cry_1), .S(mult1_un54_sum_axb_3), .Y(), 
        .FCO(mult1_un47_sum_cry_2));
    SLE \tim[3]  (.D(\mult1_un138_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[3]));
    SLE \tim[2]  (.D(\mult1_un145_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[2]));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_9  (.A(
        mult1_un68_sum_cry_8_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_8), .S(
        mult1_un75_sum_cry_9_S), .Y(), .FCO(mult1_un75_sum_cry_9));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un54_sum_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_1  (.A(\i_i[11] )
        , .B(mult1_un96_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), 
        .FCI(mult1_un103_sum_cry_0), .S(mult1_un103_sum_cry_1_S), .Y(), 
        .FCO(mult1_un103_sum_cry_1));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un145_sum_cry_10_S), .C(mult1_un145_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un152_sum_cry_10), .S(
        mult1_un152_sum_s_11_S), .Y(), .FCO());
    SLE \state[4]  (.D(N_183_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    ARI1 #( .INIT(20'h67700) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_7  (.A(VCC_net_1), 
        .B(mult1_un47_sum_cry_4), .C(mult1_un47_sum_s_5_sf), .D(
        GND_net_1), .FCI(mult1_un54_sum_cry_6), .S(
        mult1_un61_sum_axb_8), .Y(), .FCO(mult1_un54_sum_cry_7));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_3  (.A(VCC_net_1), 
        .B(mult1_un68_sum_axb_3), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_2), .S(mult1_un68_sum_cry_3_S), .Y(), .FCO(
        mult1_un68_sum_cry_3));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_9  (.A(
        mult1_un152_sum_cry_8_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_8), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_9));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_8  (.A(
        mult1_un103_sum_cry_7_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_7), .S(
        mult1_un110_sum_cry_8_S), .Y(), .FCO(mult1_un110_sum_cry_8));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un75_sum_cry_10_S), .C(mult1_un75_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un82_sum_cry_10), .S(
        mult1_un82_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_5  (.A(
        mult1_un117_sum_cry_4_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_4), .S(
        mult1_un124_sum_cry_5_S), .Y(), .FCO(mult1_un124_sum_cry_5));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_3  (.A(
        mult1_un110_sum_cry_2_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_2), .S(
        mult1_un117_sum_cry_3_S), .Y(), .FCO(mult1_un117_sum_cry_3));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un96_sum_cry_10_S), .C(mult1_un96_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un103_sum_cry_10), .S(
        mult1_un103_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un110_sum_cry_10_S), .C(mult1_un110_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un117_sum_cry_10), .S(
        mult1_un117_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_7  (.A(
        mult1_un117_sum_cry_6_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_6), .S(
        mult1_un124_sum_cry_7_S), .Y(), .FCO(mult1_un124_sum_cry_7));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_i_0[13]  (.A(
        mult1_un145_sum_s_11_S), .Y(\mult1_un145_sum_i_0[13] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_10  (.A(
        mult1_un103_sum_cry_9_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_9), .S(
        mult1_un110_sum_cry_10_S), .Y(), .FCO(mult1_un110_sum_cry_10));
    CFG1 #( .INIT(2'h1) )  \i_RNIJVQ6[12]  (.A(\i[12]_net_1 ), .Y(
        \i_i[12] ));
    SLE \i[13]  (.D(\i_s[13] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_1  (.A(\i_i[5] ), 
        .B(mult1_un138_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un145_sum_cry_0), .S(mult1_un145_sum_cry_1_S), .Y(), 
        .FCO(mult1_un145_sum_cry_1));
    ARI1 #( .INIT(20'h42200) )  \i_cry[15]  (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[14]_net_1 ), .S(\i_s[15] ), .Y(), .FCO(
        \i_cry[15]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_s_5_sf  (.A(
        \i[20]_net_1 ), .B(\i[19]_net_1 ), .C(CO2), .Y(
        mult1_un47_sum_s_5_sf));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_7  (.A(
        mult1_un131_sum_cry_6_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_6), .S(
        mult1_un138_sum_cry_7_S), .Y(), .FCO(mult1_un138_sum_cry_7));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_6  (.A(
        mult1_un152_sum_cry_5_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_5), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_6));
    SLE \tim[1]  (.D(\mult1_un152_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[1]));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_3  (.A(
        mult1_un103_sum_cry_2_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_2), .S(
        mult1_un110_sum_cry_3_S), .Y(), .FCO(mult1_un110_sum_cry_3));
    SLE \tim[5]  (.D(\mult1_un124_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[5]));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_5  (.A(
        mult1_un82_sum_cry_4_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_4), .S(
        mult1_un89_sum_cry_5_S), .Y(), .FCO(mult1_un89_sum_cry_5));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_4  (.A(
        mult1_un152_sum_cry_3_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_3), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_7  (.A(
        mult1_un68_sum_cry_6_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_6), .S(
        mult1_un75_sum_cry_7_S), .Y(), .FCO(mult1_un75_sum_cry_7));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_7  (.A(VCC_net_1), 
        .B(mult1_un54_sum_cry_6_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_6), .S(mult1_un68_sum_axb_8), .Y(), .FCO(
        mult1_un61_sum_cry_7));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un138_sum_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_8  (.A(
        mult1_un96_sum_cry_7_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_7), .S(
        mult1_un103_sum_cry_8_S), .Y(), .FCO(mult1_un103_sum_cry_8));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_10  (.A(
        mult1_un96_sum_cry_9_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_9), .S(
        mult1_un103_sum_cry_10_S), .Y(), .FCO(mult1_un103_sum_cry_10));
    SLE \i[17]  (.D(\i_s[17] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[17]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un68_sum_axb_11), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_10), .S(mult1_un68_sum_s_11_S), .Y(), .FCO()
        );
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_2  (.A(
        mult1_un152_sum_cry_1_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_1), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_2));
    SLE \tim[11]  (.D(\mult1_un82_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[11]));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_6  (.A(
        mult1_un145_sum_cry_5_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_5), .S(
        mult1_un152_sum_cry_6_S), .Y(), .FCO(mult1_un152_sum_cry_6));
    ARI1 #( .INIT(20'h42200) )  \i_cry[17]  (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[16]_net_1 ), .S(\i_s[17] ), .Y(), .FCO(
        \i_cry[17]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_6  (.A(
        mult1_un110_sum_cry_5_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_5), .S(
        mult1_un117_sum_cry_6_S), .Y(), .FCO(mult1_un117_sum_cry_6));
    CFG3 #( .INIT(8'h70) )  \state_RNO[1]  (.A(\state_ns_o2[2]_net_1 ), 
        .B(ECHO_c), .C(\state[2]_net_1 ), .Y(N_187_i_0));
    CFG4 #( .INIT(16'hCC80) )  \state_ns_o2_RNIJNK11[2]  (.A(
        \state[2]_net_1 ), .B(ECHO_c), .C(\state_ns_o2[2]_net_1 ), .D(
        \state[3]_net_1 ), .Y(N_5_i_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_8  (.A(
        mult1_un117_sum_cry_7_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_7), .S(
        mult1_un124_sum_cry_8_S), .Y(), .FCO(mult1_un124_sum_cry_8));
    SLE \i[9]  (.D(\i_s[9] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_8  (.A(
        mult1_un89_sum_cry_7_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_7), .S(
        mult1_un96_sum_cry_8_S), .Y(), .FCO(mult1_un96_sum_cry_8));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_3  (.A(
        mult1_un68_sum_cry_2_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_2), .S(
        mult1_un75_sum_cry_3_S), .Y(), .FCO(mult1_un75_sum_cry_3));
    CFG1 #( .INIT(2'h1) )  \i_RNI9GK2[9]  (.A(\i[9]_net_1 ), .Y(
        \i_i[9] ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_6  (.A(
        mult1_un68_sum_cry_5_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_5), .S(
        mult1_un75_sum_cry_6_S), .Y(), .FCO(mult1_un75_sum_cry_6));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_5  (.A(
        mult1_un131_sum_cry_4_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_4), .S(
        mult1_un138_sum_cry_5_S), .Y(), .FCO(mult1_un138_sum_cry_5));
    CFG1 #( .INIT(2'h1) )  \i_RNIL1R6[14]  (.A(\i[14]_net_1 ), .Y(
        \i_i[14] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_10  (.A(
        mult1_un82_sum_cry_9_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_9), .S(
        mult1_un89_sum_cry_10_S), .Y(), .FCO(mult1_un89_sum_cry_10));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_1  (.A(\i_i[7] ), 
        .B(mult1_un124_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un131_sum_cry_0), .S(mult1_un131_sum_cry_1_S), .Y(), 
        .FCO(mult1_un131_sum_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_10  (.A(
        mult1_un124_sum_cry_9_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_9), .S(
        mult1_un131_sum_cry_10_S), .Y(), .FCO(mult1_un131_sum_cry_10));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_8  (.A(
        mult1_un145_sum_cry_7_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_7), .S(
        mult1_un152_sum_cry_8_S), .Y(), .FCO(mult1_un152_sum_cry_8));
    CFG1 #( .INIT(2'h1) )  \i_RNI7EK2[7]  (.A(\i[7]_net_1 ), .Y(
        \i_i[7] ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_i_0[13]  (.A(
        mult1_un152_sum_s_11_S), .Y(\mult1_un152_sum_i_0[13] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_10  (.A(
        mult1_un152_sum_cry_9_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_9), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_10));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un131_sum_cry_0));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_6  (.A(
        mult1_un124_sum_cry_5_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_5), .S(
        mult1_un131_sum_cry_6_S), .Y(), .FCO(mult1_un131_sum_cry_6));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_9  (.A(
        mult1_un110_sum_cry_8_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_8), .S(
        mult1_un117_sum_cry_9_S), .Y(), .FCO(mult1_un117_sum_cry_9));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_7  (.A(
        mult1_un82_sum_cry_6_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_6), .S(
        mult1_un89_sum_cry_7_S), .Y(), .FCO(mult1_un89_sum_cry_7));
    CFG4 #( .INIT(16'h000D) )  \state_RNO[4]  (.A(
        locator_control_0_en_timer), .B(\state[0]_net_1 ), .C(
        \state_ns_i_0_0[0]_net_1 ), .D(\state[1]_net_1 ), .Y(N_183_i_0)
        );
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un138_sum_cry_10_S), .C(mult1_un138_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un145_sum_cry_10), .S(
        mult1_un145_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h40000) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_s_10  (.A(VCC_net_1), 
        .B(GND_net_1), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_9), .S(mult1_un68_sum_axb_11), .Y(), .FCO());
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_9  (.A(
        mult1_un131_sum_cry_8_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_8), .S(
        mult1_un138_sum_cry_9_S), .Y(), .FCO(mult1_un138_sum_cry_9));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_5  (.A(VCC_net_1), 
        .B(mult1_un61_sum_axb_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_4), .S(mult1_un61_sum_cry_5_S), .Y(), .FCO(
        mult1_un61_sum_cry_5));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_5  (.A(
        mult1_un89_sum_cry_4_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_4), .S(
        mult1_un96_sum_cry_5_S), .Y(), .FCO(mult1_un96_sum_cry_5));
    SLE \i_fast[19]  (.D(\i_s[19] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_fast[19]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[11]  (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[10]_net_1 ), .S(\i_s[11] ), .Y(), .FCO(
        \i_cry[11]_net_1 ));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un117_sum_cry_10_S), .C(mult1_un117_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un124_sum_cry_10), .S(
        mult1_un124_sum_s_11_S), .Y(), .FCO());
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_i_0[13]  (.A(
        mult1_un159_sum_s_11_S), .Y(\mult1_un159_sum_i_0[13] ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_6  (.A(
        mult1_un96_sum_cry_5_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_5), .S(
        mult1_un103_sum_cry_6_S), .Y(), .FCO(mult1_un103_sum_cry_6));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_6  (.A(
        mult1_un89_sum_cry_5_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_5), .S(
        mult1_un96_sum_cry_6_S), .Y(), .FCO(mult1_un96_sum_cry_6));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_6  (.A(VCC_net_1), 
        .B(mult1_un54_sum_cry_5_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_5), .S(mult1_un61_sum_cry_6_S), .Y(), .FCO(
        mult1_un61_sum_cry_6));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_9  (.A(
        mult1_un75_sum_cry_8_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_8), .S(
        mult1_un82_sum_cry_9_S), .Y(), .FCO(mult1_un82_sum_cry_9));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_10  (.A(
        mult1_un75_sum_cry_9_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_9), .S(
        mult1_un82_sum_cry_10_S), .Y(), .FCO(mult1_un82_sum_cry_10));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_10  (.A(
        mult1_un68_sum_cry_9_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_9), .S(
        mult1_un75_sum_cry_10_S), .Y(), .FCO(mult1_un75_sum_cry_10));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_6  (.A(
        mult1_un131_sum_cry_5_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_5), .S(
        mult1_un138_sum_cry_6_S), .Y(), .FCO(mult1_un138_sum_cry_6));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_10  (.A(
        mult1_un145_sum_cry_9_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_9), .S(
        mult1_un152_sum_cry_10_S), .Y(), .FCO(mult1_un152_sum_cry_10));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_5  (.A(VCC_net_1), 
        .B(mult1_un54_sum_axb_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un54_sum_cry_4), .S(mult1_un54_sum_cry_5_S), .Y(), .FCO(
        mult1_un54_sum_cry_5));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_2  (.A(
        mult1_un117_sum_cry_1_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_1), .S(
        mult1_un124_sum_cry_2_S), .Y(), .FCO(mult1_un124_sum_cry_2));
    SLE \i[15]  (.D(\i_s[15] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[15]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_2  (.A(VCC_net_1), 
        .B(mult1_un54_sum_cry_1_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_1), .S(mult1_un68_sum_axb_3), .Y(), .FCO(
        mult1_un61_sum_cry_2));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_3  (.A(
        mult1_un138_sum_cry_2_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_2), .S(
        mult1_un145_sum_cry_3_S), .Y(), .FCO(mult1_un145_sum_cry_3));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_9  (.A(
        mult1_un103_sum_cry_8_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_8), .S(
        mult1_un110_sum_cry_9_S), .Y(), .FCO(mult1_un110_sum_cry_9));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un61_sum_cry_0));
    CFG1 #( .INIT(2'h1) )  \i_RNI8FK2[8]  (.A(\i[8]_net_1 ), .Y(
        \i_i[8] ));
    SLE \tim[0]  (.D(\mult1_un159_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[0]));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_2  (.A(
        mult1_un131_sum_cry_1_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_1), .S(
        mult1_un138_sum_cry_2_S), .Y(), .FCO(mult1_un138_sum_cry_2));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_i_0[13]  (.A(
        mult1_un68_sum_s_11_S), .Y(\mult1_un68_sum_i_0[13] ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_2  (.A(
        mult1_un89_sum_cry_1_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_1), .S(
        mult1_un96_sum_cry_2_S), .Y(), .FCO(mult1_un96_sum_cry_2));
    ARI1 #( .INIT(20'h42200) )  \i_cry[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7] ), .Y(), .FCO(\i_cry[7]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_3  (.A(
        mult1_un96_sum_cry_2_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_2), .S(
        mult1_un103_sum_cry_3_S), .Y(), .FCO(mult1_un103_sum_cry_3));
    ARI1 #( .INIT(20'h42200) )  \i_cry[12]  (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[11]_net_1 ), .S(\i_s[12] ), .Y(), .FCO(
        \i_cry[12]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_6  (.A(
        mult1_un117_sum_cry_5_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_5), .S(
        mult1_un124_sum_cry_6_S), .Y(), .FCO(mult1_un124_sum_cry_6));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_8  (.A(
        mult1_un138_sum_cry_7_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_7), .S(
        mult1_un145_sum_cry_8_S), .Y(), .FCO(mult1_un145_sum_cry_8));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_i_0[13]  (.A(
        mult1_un117_sum_s_11_S), .Y(\mult1_un117_sum_i_0[13] ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[18]  (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[17]_net_1 ), .S(\i_s[18] ), .Y(), .FCO(
        \i_cry[18]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_i_0[13]  (.A(
        mult1_un82_sum_s_11_S), .Y(\mult1_un82_sum_i_0[13] ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_9  (.A(VCC_net_1), 
        .B(mult1_un54_sum_s_8_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_8), .S(mult1_un68_sum_axb_10), .Y(), .FCO(
        mult1_un61_sum_cry_9));
    ARI1 #( .INIT(20'h55555) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_1  (.A(VCC_net_1), 
        .B(\i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_0), .S(mult1_un68_sum_cry_1_S), .Y(), .FCO(
        mult1_un68_sum_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_3  (.A(
        mult1_un152_sum_cry_2_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_2), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_3));
    SLE \i[2]  (.D(\i_s[2] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    SLE \i[12]  (.D(\i_s[12] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_4  (.A(VCC_net_1), 
        .B(mult1_un61_sum_cry_3_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_3), .S(mult1_un68_sum_cry_4_S), .Y(), .FCO(
        mult1_un68_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_7  (.A(
        mult1_un75_sum_cry_6_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_6), .S(
        mult1_un82_sum_cry_7_S), .Y(), .FCO(mult1_un82_sum_cry_7));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_5  (.A(
        mult1_un110_sum_cry_4_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_4), .S(
        mult1_un117_sum_cry_5_S), .Y(), .FCO(mult1_un117_sum_cry_5));
    SLE \tim[13]  (.D(\mult1_un68_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[13]));
    ARI1 #( .INIT(20'h45500) )  \i_cry_cy[0]  (.A(VCC_net_1), .B(
        \state[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(i_cry_cy));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_6  (.A(VCC_net_1), 
        .B(mult1_un61_sum_cry_5_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_5), .S(mult1_un68_sum_cry_6_S), .Y(), .FCO(
        mult1_un68_sum_cry_6));
    SLE \i[20]  (.D(\i_s[20] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[20]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_4  (.A(VCC_net_1), 
        .B(mult1_un54_sum_cry_3_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_3), .S(mult1_un68_sum_axb_5), .Y(), .FCO(
        mult1_un61_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_4  (.A(
        mult1_un145_sum_cry_3_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_3), .S(
        mult1_un152_sum_cry_4_S), .Y(), .FCO(mult1_un152_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_2  (.A(
        mult1_un110_sum_cry_1_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_1), .S(
        mult1_un117_sum_cry_2_S), .Y(), .FCO(mult1_un117_sum_cry_2));
    CFG1 #( .INIT(2'h1) )  \i_RNIK0R6[13]  (.A(\i[13]_net_1 ), .Y(
        \i_i[13] ));
    SLE \state[3]  (.D(\state_ns[1] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \i_RNIM2R6[15]  (.A(\i[15]_net_1 ), .Y(
        \i_i[15] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_3  (.A(
        mult1_un75_sum_cry_2_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_2), .S(
        mult1_un82_sum_cry_3_S), .Y(), .FCO(mult1_un82_sum_cry_3));
    SLE \i[10]  (.D(\i_s[10] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_9  (.A(
        mult1_un82_sum_cry_8_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_8), .S(
        mult1_un89_sum_cry_9_S), .Y(), .FCO(mult1_un89_sum_cry_9));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_8  (.A(
        mult1_un124_sum_cry_7_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_7), .S(
        mult1_un131_sum_cry_8_S), .Y(), .FCO(mult1_un131_sum_cry_8));
    CFG1 #( .INIT(2'h1) )  \i_RNI6DK2[6]  (.A(\i[6]_net_1 ), .Y(
        \i_i[6] ));
    CFG1 #( .INIT(2'h1) )  \i_RNI5CK2[5]  (.A(\i[5]_net_1 ), .Y(
        \i_i[5] ));
    SLE \i[6]  (.D(\i_s[6] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[0]_net_1 ), .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_s[4] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_10  (.A(
        mult1_un117_sum_cry_9_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_9), .S(
        mult1_un124_sum_cry_10_S), .Y(), .FCO(mult1_un124_sum_cry_10));
    ARI1 #( .INIT(20'h42200) )  \i_cry[10]  (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[9]_net_1 ), .S(\i_s[10] ), .Y(), .FCO(\i_cry[10]_net_1 )
        );
    SLE \tim[12]  (.D(\mult1_un75_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[12]));
    ARI1 #( .INIT(20'h42200) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_8  (.A(
        mult1_un152_sum_cry_7_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_7), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_8));
    CFG4 #( .INIT(16'hF777) )  \state_ns_o2_0[2]  (.A(\i[18]_net_1 ), 
        .B(\i[17]_net_1 ), .C(un20_clklto16_1_net_1), .D(un20_clklt16), 
        .Y(un20_clklt20));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_8  (.A(
        mult1_un68_sum_cry_7_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_7), .S(
        mult1_un75_sum_cry_8_S), .Y(), .FCO(mult1_un75_sum_cry_8));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_3  (.A(
        mult1_un124_sum_cry_2_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_2), .S(
        mult1_un131_sum_cry_3_S), .Y(), .FCO(mult1_un131_sum_cry_3));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_5  (.A(
        mult1_un145_sum_cry_4_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_4), .S(
        mult1_un152_sum_cry_5_S), .Y(), .FCO(mult1_un152_sum_cry_5));
    SLE \i[19]  (.D(\i_s[19] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[19]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_i_0[13]  (.A(
        mult1_un103_sum_s_11_S), .Y(\mult1_un103_sum_i_0[13] ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un110_sum_cry_0));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_2  (.A(
        mult1_un145_sum_cry_1_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_1), .S(
        mult1_un152_sum_cry_2_S), .Y(), .FCO(mult1_un152_sum_cry_2));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_8  (.A(
        mult1_un82_sum_cry_7_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_7), .S(
        mult1_un89_sum_cry_8_S), .Y(), .FCO(mult1_un89_sum_cry_8));
    ARI1 #( .INIT(20'h53CAA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_1  (.A(VCC_net_1)
        , .B(mult1_un103_sum_cry_0_Y), .C(\i[10]_net_1 ), .D(
        mult1_un103_sum_s_11_S), .FCI(mult1_un110_sum_cry_0), .S(
        mult1_un110_sum_cry_1_S), .Y(), .FCO(mult1_un110_sum_cry_1));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_1  (.A(\i_i[15] ), 
        .B(mult1_un68_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un75_sum_cry_0), .S(mult1_un75_sum_cry_1_S), .Y(), .FCO(
        mult1_un75_sum_cry_1));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un152_sum_cry_10_S), .C(mult1_un152_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un159_sum_cry_10), .S(
        mult1_un159_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_6  (.A(
        mult1_un138_sum_cry_5_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_5), .S(
        mult1_un145_sum_cry_6_S), .Y(), .FCO(mult1_un145_sum_cry_6));
    SLE \tim[8]  (.D(\mult1_un103_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[8]));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_5  (.A(
        mult1_un75_sum_cry_4_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_4), .S(
        mult1_un82_sum_cry_5_S), .Y(), .FCO(mult1_un82_sum_cry_5));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_4  (.A(
        mult1_un131_sum_cry_3_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_3), .S(
        mult1_un138_sum_cry_4_S), .Y(), .FCO(mult1_un138_sum_cry_4));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un68_sum_cry_10_S), .C(mult1_un68_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un75_sum_cry_10), .S(
        mult1_un75_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_3  (.A(
        mult1_un117_sum_cry_2_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_2), .S(
        mult1_un124_sum_cry_3_S), .Y(), .FCO(mult1_un124_sum_cry_3));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un103_sum_cry_10_S), .C(mult1_un103_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un110_sum_cry_10), .S(
        mult1_un110_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_1  (.A(\i_i[6] ), 
        .B(mult1_un131_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un138_sum_cry_0), .S(mult1_un138_sum_cry_1_S), .Y(), 
        .FCO(mult1_un138_sum_cry_1));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_2  (.A(
        mult1_un75_sum_cry_1_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_1), .S(
        mult1_un82_sum_cry_2_S), .Y(), .FCO(mult1_un82_sum_cry_2));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un61_sum_cry_3  (.A(VCC_net_1), 
        .B(mult1_un61_sum_axb_3), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un61_sum_cry_2), .S(mult1_un61_sum_cry_3_S), .Y(), .FCO(
        mult1_un61_sum_cry_3));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_7  (.A(
        mult1_un124_sum_cry_6_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_6), .S(
        mult1_un131_sum_cry_7_S), .Y(), .FCO(mult1_un131_sum_cry_7));
    CFG4 #( .INIT(16'hAE0C) )  \state_ns_0[1]  (.A(
        locator_control_0_en_timer), .B(\state[3]_net_1 ), .C(ECHO_c), 
        .D(\state[4]_net_1 ), .Y(\state_ns[1] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_10  (.A(
        mult1_un110_sum_cry_9_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_9), .S(
        mult1_un117_sum_cry_10_S), .Y(), .FCO(mult1_un117_sum_cry_10));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un82_sum_cry_0));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_10  (.A(
        mult1_un131_sum_cry_9_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_9), .S(
        mult1_un138_sum_cry_10_S), .Y(), .FCO(mult1_un138_sum_cry_10));
    ARI1 #( .INIT(20'h40000) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_s_8  (.A(VCC_net_1), 
        .B(GND_net_1), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un54_sum_cry_7), .S(mult1_un54_sum_s_8_S), .Y(), .FCO());
    CFG4 #( .INIT(16'h777F) )  \state_ns_o2_4[2]  (.A(\i[8]_net_1 ), 
        .B(\i[7]_net_1 ), .C(\i[6]_net_1 ), .D(\i[5]_net_1 ), .Y(
        un20_clklt9));
    CFG4 #( .INIT(16'h0F4F) )  \state_ns_o2_2[2]  (.A(\i[11]_net_1 ), 
        .B(un20_clklt12), .C(\i[13]_net_1 ), .D(\i[12]_net_1 ), .Y(
        un20_clklt16));
    SLE new_ready (.D(\state[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_201_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(pulse_meash_0_new_ready));
    CFG3 #( .INIT(8'h01) )  un20_clklto16_1 (.A(\i[16]_net_1 ), .B(
        \i[15]_net_1 ), .C(\i[14]_net_1 ), .Y(un20_clklto16_1_net_1));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_7  (.A(
        mult1_un145_sum_cry_6_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_6), .S(
        mult1_un152_sum_cry_7_S), .Y(), .FCO(mult1_un152_sum_cry_7));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_7  (.A(
        mult1_un138_sum_cry_6_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_6), .S(
        mult1_un145_sum_cry_7_S), .Y(), .FCO(mult1_un145_sum_cry_7));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un89_sum_cry_10_S), .C(mult1_un89_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un96_sum_cry_10), .S(
        mult1_un96_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(mult1_un103_sum_cry_0_Y), .FCO(
        mult1_un103_sum_cry_0));
    SLE \i[14]  (.D(\i_s[14] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_4  (.A(
        mult1_un103_sum_cry_3_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_3), .S(
        mult1_un110_sum_cry_4_S), .Y(), .FCO(mult1_un110_sum_cry_4));
    CFG4 #( .INIT(16'h555D) )  \state_ns_o2[2]  (.A(CO2), .B(
        un20_clklt20), .C(\i[20]_net_1 ), .D(\i[19]_net_1 ), .Y(
        \state_ns_o2[2]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h69900) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_6  (.A(VCC_net_1), 
        .B(mult1_un47_sum_s_5_sf), .C(mult1_un47_sum_cry_4), .D(
        GND_net_1), .FCI(mult1_un54_sum_cry_5), .S(
        mult1_un54_sum_cry_6_S), .Y(), .FCO(mult1_un54_sum_cry_6));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_5  (.A(
        mult1_un138_sum_cry_4_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_4), .S(
        mult1_un145_sum_cry_5_S), .Y(), .FCO(mult1_un145_sum_cry_5));
    SLE \state[2]  (.D(N_5_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_10  (.A(
        mult1_un89_sum_cry_9_S), .B(mult1_un89_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un96_sum_cry_9), .S(
        mult1_un96_sum_cry_10_S), .Y(), .FCO(mult1_un96_sum_cry_10));
    SLE \state[1]  (.D(N_187_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_6  (.A(
        mult1_un75_sum_cry_5_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_5), .S(
        mult1_un82_sum_cry_6_S), .Y(), .FCO(mult1_un82_sum_cry_6));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un68_sum_cry_0));
    ARI1 #( .INIT(20'h42200) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_2  (.A(
        mult1_un138_sum_cry_1_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_1), .S(
        mult1_un145_sum_cry_2_S), .Y(), .FCO(mult1_un145_sum_cry_2));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_cry_3  (.A(
        mult1_un131_sum_cry_2_S), .B(mult1_un131_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un138_sum_cry_2), .S(
        mult1_un138_sum_cry_3_S), .Y(), .FCO(mult1_un138_sum_cry_3));
    SLE \i[5]  (.D(\i_s[5] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_6  (.A(
        mult1_un103_sum_cry_5_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_5), .S(
        mult1_un110_sum_cry_6_S), .Y(), .FCO(mult1_un110_sum_cry_6));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_7  (.A(
        mult1_un110_sum_cry_6_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_6), .S(
        mult1_un117_sum_cry_7_S), .Y(), .FCO(mult1_un117_sum_cry_7));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_2  (.A(
        mult1_un103_sum_cry_1_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_1), .S(
        mult1_un110_sum_cry_2_S), .Y(), .FCO(mult1_un110_sum_cry_2));
    SLE \i[8]  (.D(\i_s[8] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_i_0[13]  (.A(
        mult1_un96_sum_s_11_S), .Y(\mult1_un96_sum_i_0[13] ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_7  (.A(
        mult1_un96_sum_cry_6_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_6), .S(
        mult1_un103_sum_cry_7_S), .Y(), .FCO(mult1_un103_sum_cry_7));
    SLE \tim[6]  (.D(\mult1_un117_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[6]));
    ARI1 #( .INIT(20'h42200) )  \i_cry[13]  (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[12]_net_1 ), .S(\i_s[13] ), .Y(), .FCO(
        \i_cry[13]_net_1 ));
    ARI1 #( .INIT(20'h41E00) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_cry_3  (.A(VCC_net_1), 
        .B(\i_fast[19]_net_1 ), .C(\i_fast[20]_net_1 ), .D(
        \i_fast[21]_net_1 ), .FCI(mult1_un47_sum_cry_2), .S(
        mult1_un47_sum_cry_3_S), .Y(), .FCO(mult1_un47_sum_cry_3));
    SLE \tim[9]  (.D(\mult1_un96_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[9]));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_9  (.A(VCC_net_1), 
        .B(mult1_un61_sum_cry_8_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_8), .S(mult1_un68_sum_cry_9_S), .Y(), .FCO(
        mult1_un68_sum_cry_9));
    ARI1 #( .INIT(20'h53CAA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_1  (.A(VCC_net_1)
        , .B(mult1_un152_sum_cry_0_Y), .C(\i[3]_net_1 ), .D(
        mult1_un152_sum_s_11_S), .FCI(mult1_un159_sum_cry_0), .S(), .Y(
        ), .FCO(mult1_un159_sum_cry_1));
    ARI1 #( .INIT(20'h42200) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_5  (.A(VCC_net_1), 
        .B(mult1_un68_sum_axb_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_4), .S(mult1_un68_sum_cry_5_S), .Y(), .FCO(
        mult1_un68_sum_cry_5));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_3  (.A(VCC_net_1), 
        .B(mult1_un54_sum_axb_3), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un54_sum_cry_2), .S(mult1_un54_sum_cry_3_S), .Y(), .FCO(
        mult1_un54_sum_cry_3));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_5  (.A(
        mult1_un103_sum_cry_4_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_4), .S(
        mult1_un110_sum_cry_5_S), .Y(), .FCO(mult1_un110_sum_cry_5));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_9  (.A(
        mult1_un145_sum_cry_8_S), .B(mult1_un145_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un152_sum_cry_8), .S(
        mult1_un152_sum_cry_9_S), .Y(), .FCO(mult1_un152_sum_cry_9));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_9  (.A(
        mult1_un96_sum_cry_8_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_8), .S(
        mult1_un103_sum_cry_9_S), .Y(), .FCO(mult1_un103_sum_cry_9));
    SLE \tim[10]  (.D(\mult1_un89_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[10]));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_8  (.A(
        mult1_un110_sum_cry_7_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_7), .S(
        mult1_un117_sum_cry_8_S), .Y(), .FCO(mult1_un117_sum_cry_8));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_4  (.A(
        mult1_un68_sum_cry_3_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_3), .S(
        mult1_un75_sum_cry_4_S), .Y(), .FCO(mult1_un75_sum_cry_4));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un47_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(mult1_un47_sum_cry_0_Y), .FCO(
        mult1_un47_sum_cry_0));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un145_sum_cry_0));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un117_sum_cry_0));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_i_0[13]  (.A(
        mult1_un138_sum_s_11_S), .Y(\mult1_un138_sum_i_0[13] ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_5  (.A(
        mult1_un152_sum_cry_4_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_4), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_5));
    ARI1 #( .INIT(20'h42200) )  \i_cry[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[8]_net_1 ), .S(\i_s[9] ), .Y(), .FCO(\i_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un75_sum_cry_0));
    SLE \i[3]  (.D(\i_s[3] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_4  (.A(
        mult1_un117_sum_cry_3_S), .B(mult1_un117_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un124_sum_cry_3), .S(
        mult1_un124_sum_cry_4_S), .Y(), .FCO(mult1_un124_sum_cry_4));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un138_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un131_sum_cry_10_S), .C(mult1_un131_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un138_sum_cry_10), .S(
        mult1_un138_sum_s_11_S), .Y(), .FCO());
    SLE \i_fast[20]  (.D(\i_s[20] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i_fast[20]_net_1 ));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un124_sum_cry_10_S), .C(mult1_un124_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un131_sum_cry_10), .S(
        mult1_un131_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h42200) )  \i_cry[16]  (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[15]_net_1 ), .S(\i_s[16] ), .Y(), .FCO(
        \i_cry[16]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_1  (.A(\i_i[13] ), 
        .B(mult1_un82_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un89_sum_cry_0), .S(mult1_un89_sum_cry_1_S), .Y(), .FCO(
        mult1_un89_sum_cry_1));
    SLE \i_fast[21]  (.D(\i_s[21]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_5_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\i_fast[21]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_cry[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[7]_net_1 ), .S(\i_s[8] ), .Y(), .FCO(\i_cry[8]_net_1 ));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_i_0[13]  (.A(
        mult1_un75_sum_s_11_S), .Y(\mult1_un75_sum_i_0[13] ));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_2  (.A(VCC_net_1), 
        .B(mult1_un47_sum_cry_1_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un54_sum_cry_1), .S(mult1_un61_sum_axb_3), .Y(), .FCO(
        mult1_un54_sum_cry_2));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_4  (.A(
        mult1_un75_sum_cry_3_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_3), .S(
        mult1_un82_sum_cry_4_S), .Y(), .FCO(mult1_un82_sum_cry_4));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un152_sum_cry_1  (.A(\i_i[4] ), 
        .B(mult1_un145_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un152_sum_cry_0), .S(mult1_un152_sum_cry_1_S), .Y(), 
        .FCO(mult1_un152_sum_cry_1));
    ARI1 #( .INIT(20'h42200) )  \i_cry[0]  (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        i_cry_cy), .S(\i_s[0] ), .Y(), .FCO(\i_cry[0]_net_1 ));
    SLE \i[1]  (.D(\i_s[1] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    ARI1 #( .INIT(20'h533AA) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_1  (.A(VCC_net_1), 
        .B(mult1_un47_sum_cry_0_Y), .C(\i[18]_net_1 ), .D(GND_net_1), 
        .FCI(mult1_un54_sum_cry_0), .S(mult1_un54_sum_cry_1_S), .Y(), 
        .FCO(mult1_un54_sum_cry_1));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un117_sum_cry_4  (.A(
        mult1_un110_sum_cry_3_S), .B(mult1_un110_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un117_sum_cry_3), .S(
        mult1_un117_sum_cry_4_S), .Y(), .FCO(mult1_un117_sum_cry_4));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un110_sum_cry_7  (.A(
        mult1_un103_sum_cry_6_S), .B(mult1_un103_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un110_sum_cry_6), .S(
        mult1_un110_sum_cry_7_S), .Y(), .FCO(mult1_un110_sum_cry_7));
    CFG1 #( .INIT(2'h1) )  \i_RNIIUQ6[11]  (.A(\i[11]_net_1 ), .Y(
        \i_i[11] ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un145_sum_cry_9  (.A(
        mult1_un138_sum_cry_8_S), .B(mult1_un138_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un145_sum_cry_8), .S(
        mult1_un145_sum_cry_9_S), .Y(), .FCO(mult1_un145_sum_cry_9));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_2  (.A(
        mult1_un96_sum_cry_1_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_1), .S(
        mult1_un103_sum_cry_2_S), .Y(), .FCO(mult1_un103_sum_cry_2));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_6  (.A(
        mult1_un82_sum_cry_5_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_5), .S(
        mult1_un89_sum_cry_6_S), .Y(), .FCO(mult1_un89_sum_cry_6));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un159_sum_cry_7  (.A(
        mult1_un152_sum_cry_6_S), .B(mult1_un152_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un159_sum_cry_6), .S(), 
        .Y(), .FCO(mult1_un159_sum_cry_7));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_0  (.A(VCC_net_1), 
        .B(\i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un96_sum_cry_0));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un75_sum_cry_2  (.A(
        mult1_un68_sum_cry_1_S), .B(mult1_un68_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un75_sum_cry_1), .S(
        mult1_un75_sum_cry_2_S), .Y(), .FCO(mult1_un75_sum_cry_2));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_9  (.A(
        mult1_un124_sum_cry_8_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_8), .S(
        mult1_un131_sum_cry_9_S), .Y(), .FCO(mult1_un131_sum_cry_9));
    ARI1 #( .INIT(20'h49900) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_s_11  (.A(VCC_net_1), 
        .B(mult1_un82_sum_cry_10_S), .C(mult1_un82_sum_s_11_S), .D(
        GND_net_1), .FCI(mult1_un89_sum_cry_10), .S(
        mult1_un89_sum_s_11_S), .Y(), .FCO());
    ARI1 #( .INIT(20'h42200) )  \i_cry[19]  (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(\state[3]_net_1 ), .D(GND_net_1), .FCI(
        \i_cry[18]_net_1 ), .S(\i_s[19] ), .Y(), .FCO(
        \i_cry[19]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un82_sum_cry_8  (.A(
        mult1_un75_sum_cry_7_S), .B(mult1_un75_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un82_sum_cry_7), .S(
        mult1_un82_sum_cry_8_S), .Y(), .FCO(mult1_un82_sum_cry_8));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un103_sum_cry_5  (.A(
        mult1_un96_sum_cry_4_S), .B(mult1_un96_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un103_sum_cry_4), .S(
        mult1_un103_sum_cry_5_S), .Y(), .FCO(mult1_un103_sum_cry_5));
    SLE \i[18]  (.D(\i_s[18] ), .CLK(FCCC_0_GL0), .EN(N_5_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[18]_net_1 ));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_cry_2  (.A(
        mult1_un124_sum_cry_1_S), .B(mult1_un124_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un131_sum_cry_1), .S(
        mult1_un131_sum_cry_2_S), .Y(), .FCO(mult1_un131_sum_cry_2));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un124_sum_cry_0  (.A(VCC_net_1)
        , .B(\i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(mult1_un124_sum_cry_0));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un54_sum_cry_4  (.A(VCC_net_1), 
        .B(mult1_un47_sum_cry_3_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un54_sum_cry_3), .S(mult1_un61_sum_axb_5), .Y(), .FCO(
        mult1_un54_sum_cry_4));
    ARI1 #( .INIT(20'h5AA55) )  
        \un5_tim.if_generate_plus.mult1_un96_sum_cry_1  (.A(\i_i[12] ), 
        .B(mult1_un89_sum_s_11_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un96_sum_cry_0), .S(mult1_un96_sum_cry_1_S), .Y(), .FCO(
        mult1_un96_sum_cry_1));
    ARI1 #( .INIT(20'h5AAAA) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_8  (.A(VCC_net_1), 
        .B(mult1_un68_sum_axb_8), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_7), .S(mult1_un68_sum_cry_8_S), .Y(), .FCO(
        mult1_un68_sum_cry_8));
    ARI1 #( .INIT(20'h65500) )  
        \un5_tim.if_generate_plus.mult1_un68_sum_cry_7  (.A(VCC_net_1), 
        .B(mult1_un61_sum_cry_6_S), .C(GND_net_1), .D(GND_net_1), .FCI(
        mult1_un68_sum_cry_6), .S(mult1_un68_sum_cry_7_S), .Y(), .FCO(
        mult1_un68_sum_cry_7));
    CFG1 #( .INIT(2'h1) )  
        \un5_tim.if_generate_plus.mult1_un131_sum_i_0[13]  (.A(
        mult1_un131_sum_s_11_S), .Y(\mult1_un131_sum_i_0[13] ));
    CFG2 #( .INIT(4'hE) )  new_ready_RNO (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(N_201_i_0));
    ARI1 #( .INIT(20'h555AA) )  
        \un5_tim.if_generate_plus.mult1_un89_sum_cry_4  (.A(
        mult1_un82_sum_cry_3_S), .B(mult1_un82_sum_s_11_S), .C(
        GND_net_1), .D(GND_net_1), .FCI(mult1_un89_sum_cry_3), .S(
        mult1_un89_sum_cry_4_S), .Y(), .FCO(mult1_un89_sum_cry_4));
    SLE \tim[7]  (.D(\mult1_un110_sum_i_0[13] ), .CLK(FCCC_0_GL0), .EN(
        \state[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pulse_meash_0_tim[7]));
    
endmodule


module locator_control(
       BT_module_0_data_buf,
       locator_control_0_angle1,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       un46_clk_0,
       un46_clk_1,
       un46_clk_2,
       un46_clk_3,
       TRIG_c,
       locator_control_0_en_timer,
       pulse_meash_0_new_ready,
       N_234_0
    );
input  [7:0] BT_module_0_data_buf;
output [3:0] locator_control_0_angle1;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
output un46_clk_0;
output un46_clk_1;
output un46_clk_2;
output un46_clk_3;
output TRIG_c;
output locator_control_0_en_timer;
input  pulse_meash_0_new_ready;
output N_234_0;

    wire \i[26]_net_1 , VCC_net_1, \i_4_i_i_a3[26]_net_1 , N_243_i_0, 
        GND_net_1, \i[27]_net_1 , \i_4_i_i_a3[27]_net_1 , 
        \i[28]_net_1 , \i_4_i_i_a3[28]_net_1 , \i[29]_net_1 , 
        \i_4_i_i_a3[29]_net_1 , \i[30]_net_1 , \i_4_i_i_a3[30]_net_1 , 
        \st_angle[0]_net_1 , fn_angle_0_sqmuxa_net_1, 
        \st_angle[1]_net_1 , \st_angle[2]_net_1 , \st_angle[3]_net_1 , 
        un38_clk_0, un38_clk_1, un38_clk_2, un38_clk_3, \i[11]_net_1 , 
        N_458, \i[12]_net_1 , N_459, \i[13]_net_1 , N_460, 
        \i[14]_net_1 , N_461, \i[15]_net_1 , N_462, \i[16]_net_1 , 
        N_463, \i[17]_net_1 , N_464, \i[18]_net_1 , N_465, 
        \i[19]_net_1 , N_466, \i[20]_net_1 , N_467, \i[21]_net_1 , 
        \i_4_i_i_a3[21]_net_1 , \i[22]_net_1 , \i_4_i_i_a3[22]_net_1 , 
        \i[23]_net_1 , \i_4_i_i_a3[23]_net_1 , \i[24]_net_1 , 
        \i_4_i_i_a3[24]_net_1 , \i[25]_net_1 , \i_4_i_i_a3[25]_net_1 , 
        \i[0]_net_1 , N_230, \i[1]_net_1 , N_231, \i[2]_net_1 , N_232, 
        \i[3]_net_1 , N_233, \i[4]_net_1 , N_234, \i[5]_net_1 , N_235, 
        \i[6]_net_1 , N_455, \i[7]_net_1 , N_456, \i[8]_net_1 , N_457, 
        \i[9]_net_1 , N_241, \i[10]_net_1 , N_242, \state[4]_net_1 , 
        over_net_1, over_1_sqmuxa, un1_angle_0_sqmuxa_0_0_net_1, 
        \state[8]_net_1 , un1_state_8_i_0, dir_net_1, 
        cr_angle_1_sqmuxa, un1_cr_angle_1_sqmuxa_0_0_net_1, 
        \state[6]_net_1 , N_244_i_0, \state[5]_net_1 , 
        \state[3]_net_1 , \state_ns[8]_net_1 , \state[2]_net_1 , 
        N_211_i_0, \state[1]_net_1 , \state[0]_net_1 , \state_ns[11] , 
        \state[11]_net_1 , N_195_i_0, \state[10]_net_1 , 
        \state[9]_net_1 , N_201_i_0, \state[7]_net_1 , \state_ns[4] , 
        N_204_i_0, \cr_angle_s[0] , \cr_angle_s[1] , \cr_angle_s[2] , 
        \cr_angle_s[3] , un46_clk_4, \cr_angle_s[4] , un46_clk_5, 
        \cr_angle_s[5] , un46_clk_6, \cr_angle_s[6] , un46_clk_7, 
        \cr_angle_s[7] , un46_clk_8, \cr_angle_s[8] , un46_clk_9, 
        \cr_angle_s[9] , un46_clk_10, \cr_angle_s[10] , un46_clk_11, 
        \cr_angle_s[11] , un46_clk_12, \cr_angle_s[12] , un46_clk_13, 
        \cr_angle_s[13] , un46_clk_14, \cr_angle_s[14] , un46_clk_15, 
        \cr_angle_s[15] , un46_clk_16, \cr_angle_s[16] , un46_clk_17, 
        \cr_angle_s[17] , un46_clk_18, \cr_angle_s[18] , un46_clk_19, 
        \cr_angle_s[19] , un46_clk_20, \cr_angle_s[20] , un46_clk_21, 
        \cr_angle_s[21] , un46_clk_22, \cr_angle_s[22] , un46_clk_23, 
        \cr_angle_s[23] , un46_clk_24, \cr_angle_s[24] , un46_clk_25, 
        \cr_angle_s[25] , un46_clk_26, \cr_angle_s[26] , un46_clk_27, 
        \cr_angle_s[27] , un46_clk_28, \cr_angle_s[28] , un46_clk_29, 
        \cr_angle_s[29] , un46_clk_30, \cr_angle_s[30] , 
        cr_angle_lcry_cy, un38_clk_cry_30_net_1, N_229, N_291, 
        cr_angle, un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y, N_191_i_0_0, 
        N_451_i_0, \cr_angle_cry[0] , \cr_angle_lxu;_0[0] , 
        \cr_angle_qxu[0]_net_1 , \cr_angle_cry[1] , N_191_i_0, 
        \cr_angle_cry[2] , \cr_angle_cry[3] , \cr_angle_cry[4] , 
        \cr_angle_cry[5] , \cr_angle_cry[6] , \cr_angle_cry[7] , 
        \cr_angle_cry[8] , \cr_angle_cry[9] , \cr_angle_cry[10] , 
        \cr_angle_cry[11] , \cr_angle_cry[12] , \cr_angle_cry[13] , 
        \cr_angle_cry[14] , \cr_angle_cry[15] , \cr_angle_cry[16] , 
        \cr_angle_cry[17] , \cr_angle_cry[18] , \cr_angle_cry[19] , 
        \cr_angle_cry[20] , \cr_angle_cry[21] , \cr_angle_cry[22] , 
        \cr_angle_cry[23] , \cr_angle_cry[24] , \cr_angle_cry[25] , 
        \cr_angle_cry[26] , \cr_angle_cry[27] , \cr_angle_cry[28] , 
        \cr_angle_cry[29] , un46_clk_cry_0_net_1, un46_clk_cry_1_net_1, 
        un46_clk_cry_2_net_1, un46_clk_cry_3_net_1, 
        un46_clk_cry_4_net_1, un46_clk_cry_5_net_1, 
        un46_clk_cry_6_net_1, un46_clk_cry_7_net_1, 
        un46_clk_cry_8_net_1, un46_clk_cry_9_net_1, 
        un46_clk_cry_10_net_1, un46_clk_cry_11_net_1, 
        un46_clk_cry_12_net_1, un46_clk_cry_13_net_1, 
        un46_clk_cry_14_net_1, un46_clk_cry_15_net_1, 
        un46_clk_cry_16_net_1, un46_clk_cry_17_net_1, 
        un46_clk_cry_18_net_1, un46_clk_cry_19_net_1, 
        un46_clk_cry_20_net_1, un46_clk_cry_21_net_1, 
        un46_clk_cry_22_net_1, un46_clk_cry_23_net_1, 
        un46_clk_cry_24_net_1, un46_clk_cry_25_net_1, 
        un46_clk_cry_26_net_1, un46_clk_cry_27_net_1, 
        un46_clk_cry_28_net_1, un46_clk_cry_29_net_1, 
        un46_clk_cry_30_net_1, un38_clk_cry_0_net_1, 
        un38_clk_cry_1_net_1, un38_clk_cry_2_net_1, 
        un38_clk_cry_3_net_1, un38_clk_cry_4_net_1, 
        un38_clk_cry_5_net_1, un38_clk_cry_6_net_1, 
        un38_clk_cry_7_net_1, un38_clk_cry_8_net_1, 
        un38_clk_cry_9_net_1, un38_clk_cry_10_net_1, 
        un38_clk_cry_11_net_1, un38_clk_cry_12_net_1, 
        un38_clk_cry_13_net_1, un38_clk_cry_14_net_1, 
        un38_clk_cry_15_net_1, un38_clk_cry_16_net_1, 
        un38_clk_cry_17_net_1, un38_clk_cry_18_net_1, 
        un38_clk_cry_19_net_1, un38_clk_cry_20_net_1, 
        un38_clk_cry_21_net_1, un38_clk_cry_22_net_1, 
        un38_clk_cry_23_net_1, un38_clk_cry_24_net_1, 
        un38_clk_cry_25_net_1, un38_clk_cry_26_net_1, 
        un38_clk_cry_27_net_1, un38_clk_cry_28_net_1, 
        un38_clk_cry_29_net_1, un1_i_s_1_322_FCO, un1_i_cry_1_net_1, 
        un1_i_cry_1_S, un1_i_cry_2_net_1, un1_i_cry_2_S, 
        un1_i_cry_3_net_1, un1_i_cry_3_S, un1_i_cry_4_net_1, 
        un1_i_cry_4_S, un1_i_cry_5_net_1, un1_i_cry_5_S, 
        un1_i_cry_6_net_1, un1_i_cry_6_S, un1_i_cry_7_net_1, 
        un1_i_cry_7_S, un1_i_cry_8_net_1, un31_clklto8, 
        un1_i_cry_9_net_1, un1_i_cry_9_S, un1_i_cry_10_net_1, 
        un1_i_cry_10_S, un1_i_cry_11_net_1, un1_i_cry_11_S, 
        un1_i_cry_12_net_1, un1_i_cry_12_S, un1_i_cry_13_net_1, 
        un1_i_cry_13_S, un1_i_cry_14_net_1, un1_i_cry_14_S, 
        un1_i_cry_15_net_1, un1_i_cry_15_S, un1_i_cry_16_net_1, 
        un1_i_cry_16_S, un1_i_cry_17_net_1, un31_clklto17, 
        un1_i_cry_18_net_1, un1_i_cry_18_S, un1_i_cry_19_net_1, 
        un1_i_cry_19_S, un1_i_cry_20_net_1, un31_clklto20, 
        un1_i_cry_21_net_1, un31_clklto21, un1_i_cry_22_net_1, 
        un1_i_cry_22_S, un1_i_cry_23_net_1, un1_i_cry_23_S, 
        un1_i_cry_24_net_1, un1_i_cry_24_S, un1_i_cry_25_net_1, 
        un1_i_cry_25_S, un1_i_cry_26_net_1, un1_i_cry_26_S, 
        un1_i_cry_27_net_1, un1_i_cry_27_S, un1_i_cry_28_net_1, 
        un1_i_cry_28_S, un1_i_s_30_S, un1_i_cry_29_net_1, 
        un1_i_cry_29_S, \cr_angle_lxu;[0] , N_503, N_449_5, 
        \state_ns_a2_0_0_a3_0_6[8]_net_1 , 
        \state_ns_a2_0_0_a3_0_5[8]_net_1 , 
        un1_state_8_0_0_a3_10_3_net_1, un1_state_8_0_0_a3_10_2_net_1, 
        \state_ns_a2_0_0_a2_0_6[8]_net_1 , 
        \state_ns_a2_0_0_a2_0_5[8]_net_1 , un1_state_8_0_0_o2_2_net_1, 
        \state_ns_a2_0_a2_5[4]_net_1 , \state_ns_a2_0_a2_4[4]_net_1 , 
        \state_ns_i_0_0_a2_4_1[3]_net_1 , N_316, N_59, N_482, 
        \state_ns_a2_0_0_a3_0_7[8]_net_1 , un1_state_8_0_0_o2_net_1, 
        N_311, N_258, N_484, N_109, N_192, N_112, N_449_9, N_446, 
        N_116, N_114, N_117, N_452_1, N_118, N_120, N_491, N_481;
    
    CFG2 #( .INIT(4'h8) )  un1_angle_0_sqmuxa_0_0_a3 (.A(over_net_1), 
        .B(\state[1]_net_1 ), .Y(N_195_i_0));
    SLE \cr_angle[21]  (.D(\cr_angle_s[21] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_21));
    SLE \state[0]  (.D(\state_ns[11] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    SLE \cr_angle[8]  (.D(\cr_angle_s[8] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_8));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_9 (.A(VCC_net_1), .B(
        un46_clk_9), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_8_net_1), .S(), .Y(), .FCO(un46_clk_cry_9_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIDIPI21[15]  (.A(N_191_i_0)
        , .B(un46_clk_15), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[14] ), .S(\cr_angle_s[15] ), .Y(), .FCO(
        \cr_angle_cry[15] ));
    ARI1 #( .INIT(20'h5CCAA) )  \cr_angle_qxu_RNIL3NT3[0]  (.A(
        VCC_net_1), .B(\cr_angle_lxu;_0[0] ), .C(
        \cr_angle_qxu[0]_net_1 ), .D(GND_net_1), .FCI(cr_angle), .S(
        \cr_angle_s[0] ), .Y(), .FCO(\cr_angle_cry[0] ));
    SLE \i[7]  (.D(N_456), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_29 (.A(VCC_net_1), .B(
        un46_clk_29), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_28_net_1), .S(), .Y(), .FCO(un46_clk_cry_29_net_1)
        );
    SLE \angle1[2]  (.D(un46_clk_2), .CLK(FCCC_0_GL0), .EN(
        \state[4]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        locator_control_0_angle1[2]));
    SLE \i[16]  (.D(N_463), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[16]_net_1 ));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIG836B1[21]  (.A(N_191_i_0)
        , .B(un46_clk_21), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[20] ), .S(\cr_angle_s[21] ), .Y(), .FCO(
        \cr_angle_cry[21] ));
    CFG3 #( .INIT(8'hAE) )  \state_ns_o2_0_0_o3[11]  (.A(
        \state[9]_net_1 ), .B(\state[1]_net_1 ), .C(over_net_1), .Y(
        N_234_0));
    SLE \fn_angle[1]  (.D(BT_module_0_data_buf[5]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un38_clk_1));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_18 (.A(VCC_net_1), .B(
        un46_clk_18), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_17_net_1), .S(), .Y(), .FCO(un38_clk_cry_18_net_1)
        );
    SLE \cr_angle[23]  (.D(\cr_angle_s[23] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_23));
    SLE \i[21]  (.D(\i_4_i_i_a3[21]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[21]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[26]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_26_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[26]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[18]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_18_S), .C(N_446), .D(N_481), .Y(N_465));
    CFG2 #( .INIT(4'h4) )  cr_angle_1_sqmuxa_0_a3_0_a3 (.A(
        un38_clk_cry_30_net_1), .B(N_291), .Y(cr_angle_1_sqmuxa));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_26 (.A(VCC_net_1), .B(
        un46_clk_26), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_25_net_1), .S(), .Y(), .FCO(un46_clk_cry_26_net_1)
        );
    ARI1 #( .INIT(20'h5AA55) )  un38_clk_cry_0 (.A(un38_clk_0), .B(
        un46_clk_0), .C(GND_net_1), .D(GND_net_1), .FCI(GND_net_1), .S(
        ), .Y(), .FCO(un38_clk_cry_0_net_1));
    SLE \state[10]  (.D(\state[11]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[10]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[2]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_2_S), .C(N_446), .D(N_481), .Y(N_232));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI79EDR[10]  (.A(N_191_i_0), 
        .B(un46_clk_10), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[9] ), .S(\cr_angle_s[10] ), .Y(), .FCO(
        \cr_angle_cry[10] ));
    SLE \i[0]  (.D(N_230), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_a2_0_0_a3_0_6[8]  (.A(
        un1_i_cry_5_S), .B(un31_clklto8), .C(un1_i_cry_1_S), .D(
        un1_i_cry_4_S), .Y(\state_ns_a2_0_0_a3_0_6[8]_net_1 ));
    SLE \i[11]  (.D(N_458), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    ARI1 #( .INIT(20'h46A00) )  \cr_angle_RNO[30]  (.A(VCC_net_1), .B(
        N_191_i_0), .C(un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y), .D(
        un46_clk_30), .FCI(\cr_angle_cry[29] ), .S(\cr_angle_s[30] ), 
        .Y(), .FCO());
    ARI1 #( .INIT(20'h5AA55) )  un46_clk_cry_3 (.A(un46_clk_3), .B(
        \st_angle[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_2_net_1), .S(), .Y(), .FCO(un46_clk_cry_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_s_30 (.A(VCC_net_1), .B(
        \i[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_29_net_1), .S(un1_i_s_30_S), .Y(), .FCO());
    SLE \state[6]  (.D(N_204_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[6]_net_1 ));
    CFG4 #( .INIT(16'hDFFF) )  \state_ns_a2_0_0_o2_2[8]  (.A(
        un1_i_cry_16_S), .B(N_484), .C(un1_i_cry_14_S), .D(
        un1_i_cry_15_S), .Y(N_112));
    SLE dir (.D(cr_angle_1_sqmuxa), .CLK(FCCC_0_GL0), .EN(
        un1_cr_angle_1_sqmuxa_0_0_net_1), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(dir_net_1));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_11 (.A(VCC_net_1), .B(
        un46_clk_11), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_10_net_1), .S(), .Y(), .FCO(un46_clk_cry_11_net_1)
        );
    SLE \st_angle[2]  (.D(BT_module_0_data_buf[2]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \st_angle[2]_net_1 ));
    SLE \angle1[1]  (.D(un46_clk_1), .CLK(FCCC_0_GL0), .EN(
        \state[4]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        locator_control_0_angle1[1]));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIE0NTG1[25]  (.A(N_191_i_0)
        , .B(un46_clk_25), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[24] ), .S(\cr_angle_s[25] ), .Y(), .FCO(
        \cr_angle_cry[25] ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_21 (.A(VCC_net_1), .B(
        un46_clk_21), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_20_net_1), .S(), .Y(), .FCO(un38_clk_cry_21_net_1)
        );
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_19 (.A(VCC_net_1), .B(
        un46_clk_19), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_18_net_1), .S(), .Y(), .FCO(un38_clk_cry_19_net_1)
        );
    CFG2 #( .INIT(4'h7) )  \state_RNILFEF[10]  (.A(\state[10]_net_1 ), 
        .B(FCCC_0_LOCK), .Y(N_451_i_0));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[23]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_23_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[23]_net_1 ));
    CFG4 #( .INIT(16'hB8F0) )  \cr_angle_lxu[0]  (.A(
        \st_angle[0]_net_1 ), .B(FCCC_0_LOCK), .C(un46_clk_0), .D(
        \state[10]_net_1 ), .Y(\cr_angle_lxu;[0] ));
    ARI1 #( .INIT(20'h5AA55) )  un46_clk_cry_0 (.A(un46_clk_0), .B(
        \st_angle[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(), .FCO(un46_clk_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_23 (.A(VCC_net_1), .B(
        \i[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_22_net_1), .S(un1_i_cry_23_S), .Y(), .FCO(
        un1_i_cry_23_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIU40KC1[22]  (.A(N_191_i_0)
        , .B(un46_clk_22), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[21] ), .S(\cr_angle_s[22] ), .Y(), .FCO(
        \cr_angle_cry[22] ));
    CFG4 #( .INIT(16'h0F4F) )  \state_ns_i_0_0_o2_5[3]  (.A(
        \i[2]_net_1 ), .B(\state_ns_i_0_0_a2_4_1[3]_net_1 ), .C(
        \i[5]_net_1 ), .D(\i[3]_net_1 ), .Y(N_109));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[5]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_5_S), .C(N_446), .D(N_481), .Y(N_235));
    SLE \cr_angle[2]  (.D(\cr_angle_s[2] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_2));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI75E7L1[28]  (.A(N_191_i_0)
        , .B(un46_clk_28), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[27] ), .S(\cr_angle_s[28] ), .Y(), .FCO(
        \cr_angle_cry[28] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_21 (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_20_net_1), .S(un31_clklto21), .Y(), .FCO(
        un1_i_cry_21_net_1));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[15]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_15_S), .C(N_446), .D(N_481), .Y(N_462));
    SLE \cr_angle[14]  (.D(\cr_angle_s[14] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_14));
    CFG2 #( .INIT(4'h2) )  un1_cr_angle_1_sqmuxa_0_0_a2 (.A(
        \state[2]_net_1 ), .B(dir_net_1), .Y(N_291));
    CFG3 #( .INIT(8'h75) )  \state_ns_i_0_0_o2_3[3]  (.A(\i[10]_net_1 )
        , .B(\i[9]_net_1 ), .C(N_116), .Y(N_117));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_20 (.A(VCC_net_1), .B(
        un46_clk_20), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_19_net_1), .S(), .Y(), .FCO(un38_clk_cry_20_net_1)
        );
    SLE \cr_angle[6]  (.D(\cr_angle_s[6] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_6));
    SLE \state[4]  (.D(\state[5]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[24]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_24_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[24]_net_1 ));
    CFG2 #( .INIT(4'h1) )  en_sonar_RNO (.A(N_446), .B(N_503), .Y(
        un1_state_8_i_0));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[8]  (.A(\state[3]_net_1 ), 
        .B(un31_clklto8), .C(N_446), .D(N_481), .Y(N_457));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[29]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_29_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[29]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_30 (.A(VCC_net_1), .B(
        un46_clk_30), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_29_net_1), .S(), .Y(), .FCO(un38_clk_cry_30_net_1)
        );
    CFG4 #( .INIT(16'hF777) )  \state_ns_i_0_0_o2_0[3]  (.A(
        \i[17]_net_1 ), .B(\i[18]_net_1 ), .C(N_118), .D(N_59), .Y(
        N_120));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h01) )  \state_ns_a2_0_0_a3_0_5[8]  (.A(
        un1_i_cry_3_S), .B(un31_clklto20), .C(un1_i_cry_2_S), .Y(
        \state_ns_a2_0_0_a3_0_5[8]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_23 (.A(VCC_net_1), .B(
        un46_clk_23), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_22_net_1), .S(), .Y(), .FCO(un46_clk_cry_23_net_1)
        );
    SLE \state[7]  (.D(\state_ns[4] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[7]_net_1 ));
    SLE \i[23]  (.D(\i_4_i_i_a3[23]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[23]_net_1 ));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIEO1NV[13]  (.A(N_191_i_0), 
        .B(un46_clk_13), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[12] ), .S(\cr_angle_s[13] ), .Y(), .FCO(
        \cr_angle_cry[13] ));
    SLE \cr_angle[18]  (.D(\cr_angle_s[18] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_18));
    SLE \cr_angle[27]  (.D(\cr_angle_s[27] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_27));
    SLE \state[5]  (.D(\state[6]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[5]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_a2_0_0_a2_0_6[8]  (.A(
        un1_i_cry_25_S), .B(un1_i_cry_26_S), .C(un1_i_cry_27_S), .D(
        un1_i_cry_28_S), .Y(\state_ns_a2_0_0_a2_0_6[8]_net_1 ));
    SLE \cr_angle[22]  (.D(\cr_angle_s[22] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_22));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_29 (.A(VCC_net_1), .B(
        \i[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_28_net_1), .S(un1_i_cry_29_S), .Y(), .FCO(
        un1_i_cry_29_net_1));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[30]  (.A(\state[3]_net_1 ), 
        .B(un1_i_s_30_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[30]_net_1 ));
    SLE \cr_angle[29]  (.D(\cr_angle_s[29] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_29));
    SLE \i[13]  (.D(N_460), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_4 (.A(VCC_net_1), .B(
        un46_clk_4), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_3_net_1), .S(), .Y(), .FCO(un38_clk_cry_4_net_1));
    SLE \i[27]  (.D(\i_4_i_i_a3[27]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[27]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un46_clk_cry_1 (.A(un46_clk_1), .B(
        \st_angle[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_0_net_1), .S(), .Y(), .FCO(un46_clk_cry_1_net_1));
    CFG4 #( .INIT(16'h8000) )  un1_state_8_0_0_a3 (.A(N_449_5), .B(
        \state[7]_net_1 ), .C(N_449_9), .D(un1_state_8_0_0_o2_net_1), 
        .Y(N_446));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_12 (.A(VCC_net_1), .B(
        un46_clk_12), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_11_net_1), .S(), .Y(), .FCO(un46_clk_cry_12_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[28]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_28_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[28]_net_1 ));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNISGIVP[9]  (.A(N_191_i_0), 
        .B(un46_clk_9), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[8] ), .S(\cr_angle_s[9] ), .Y(), .FCO(
        \cr_angle_cry[9] ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_17 (.A(VCC_net_1), .B(
        un46_clk_17), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_16_net_1), .S(), .Y(), .FCO(un38_clk_cry_17_net_1)
        );
    ARI1 #( .INIT(20'h51BE4) )  \st_angle_RNIPT91H[3]  (.A(N_191_i_0), 
        .B(un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y), .C(
        \st_angle[3]_net_1 ), .D(un46_clk_3), .FCI(\cr_angle_cry[2] ), 
        .S(\cr_angle_s[3] ), .Y(), .FCO(\cr_angle_cry[3] ));
    SLE \i[17]  (.D(N_464), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[17]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \state_ns_i_0_0_a2_4_1[3]  (.A(
        \i[4]_net_1 ), .B(\i[0]_net_1 ), .C(\i[1]_net_1 ), .Y(
        \state_ns_i_0_0_a2_4_1[3]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_6 (.A(VCC_net_1), .B(
        un46_clk_6), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_5_net_1), .S(), .Y(), .FCO(un46_clk_cry_6_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_7 (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_6_net_1), .S(un1_i_cry_7_S), .Y(), .FCO(
        un1_i_cry_7_net_1));
    ARI1 #( .INIT(20'h51BE4) )  \st_angle_RNIVKI98[1]  (.A(N_191_i_0), 
        .B(un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y), .C(
        \st_angle[1]_net_1 ), .D(un46_clk_1), .FCI(\cr_angle_cry[0] ), 
        .S(\cr_angle_s[1] ), .Y(), .FCO(\cr_angle_cry[1] ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_8 (.A(VCC_net_1), .B(
        un46_clk_8), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_7_net_1), .S(), .Y(), .FCO(un46_clk_cry_8_net_1));
    CFG4 #( .INIT(16'hBFFF) )  un38_clk_cry_30_RNILS9U (.A(dir_net_1), 
        .B(FCCC_0_LOCK), .C(un38_clk_cry_30_net_1), .D(
        \state[2]_net_1 ), .Y(N_191_i_0));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_4 (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_3_net_1), .S(un1_i_cry_4_S), .Y(), .FCO(
        un1_i_cry_4_net_1));
    CFG2 #( .INIT(4'h8) )  fn_angle_0_sqmuxa (.A(FCCC_0_LOCK), .B(
        \state[11]_net_1 ), .Y(fn_angle_0_sqmuxa_net_1));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_12 (.A(VCC_net_1), .B(
        un46_clk_12), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_11_net_1), .S(), .Y(), .FCO(un38_clk_cry_12_net_1)
        );
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNITKT411[14]  (.A(N_191_i_0)
        , .B(un46_clk_14), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[13] ), .S(\cr_angle_s[14] ), .Y(), .FCO(
        \cr_angle_cry[14] ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_21 (.A(VCC_net_1), .B(
        un46_clk_21), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_20_net_1), .S(), .Y(), .FCO(un46_clk_cry_21_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[1]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_1_S), .C(N_446), .D(N_481), .Y(N_231));
    ARI1 #( .INIT(20'h5AA55) )  un38_clk_cry_2 (.A(un38_clk_2), .B(
        un46_clk_2), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_1_net_1), .S(), .Y(), .FCO(un38_clk_cry_2_net_1));
    SLE \i[9]  (.D(N_241), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_state_8_0_0_a3_10 (.A(
        un1_state_8_0_0_a3_10_2_net_1), .B(N_258), .C(N_59), .D(
        un1_state_8_0_0_a3_10_3_net_1), .Y(N_449_9));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_8 (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_7_net_1), .S(un31_clklto8), .Y(), .FCO(
        un1_i_cry_8_net_1));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_30 (.A(VCC_net_1), .B(
        un46_clk_30), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_29_net_1), .S(), .Y(), .FCO(un46_clk_cry_30_net_1)
        );
    ARI1 #( .INIT(20'h5AA55) )  un38_clk_cry_3 (.A(un38_clk_3), .B(
        un46_clk_3), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_2_net_1), .S(), .Y(), .FCO(un38_clk_cry_3_net_1));
    CFG3 #( .INIT(8'h01) )  \state_ns_a2_0_a2_4[4]  (.A(\i[30]_net_1 ), 
        .B(\i[27]_net_1 ), .C(\i[23]_net_1 ), .Y(
        \state_ns_a2_0_a2_4[4]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h070F) )  un46_clk_cry_30_RNIDVNA1 (.A(dir_net_1), 
        .B(\state[2]_net_1 ), .C(\state[10]_net_1 ), .D(
        un46_clk_cry_30_net_1), .Y(N_229));
    SLE \cr_angle[10]  (.D(\cr_angle_s[10] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_10));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_12 (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_11_net_1), .S(un1_i_cry_12_S), .Y(), .FCO(
        un1_i_cry_12_net_1));
    CFG4 #( .INIT(16'hF070) )  \state_ns_a2_0_0_a2_10[8]  (.A(
        un1_i_cry_10_S), .B(un1_i_cry_9_S), .C(N_316), .D(N_482), .Y(
        N_484));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[25]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_25_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[25]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_a2_0_a2_5[4]  (.A(
        \i[29]_net_1 ), .B(\i[28]_net_1 ), .C(\i[25]_net_1 ), .D(
        \i[22]_net_1 ), .Y(\state_ns_a2_0_a2_5[4]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_15 (.A(VCC_net_1), .B(
        un46_clk_15), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_14_net_1), .S(), .Y(), .FCO(un38_clk_cry_15_net_1)
        );
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_24 (.A(VCC_net_1), .B(
        un46_clk_24), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_23_net_1), .S(), .Y(), .FCO(un38_clk_cry_24_net_1)
        );
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_17 (.A(VCC_net_1), .B(
        un46_clk_17), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_16_net_1), .S(), .Y(), .FCO(un46_clk_cry_17_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_5 (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_4_net_1), .S(un1_i_cry_5_S), .Y(), .FCO(
        un1_i_cry_5_net_1));
    CFG3 #( .INIT(8'h01) )  \state_ns_a2_0_0_a2_1[8]  (.A(
        un1_i_cry_11_S), .B(un1_i_cry_12_S), .C(un1_i_cry_13_S), .Y(
        N_316));
    CFG4 #( .INIT(16'h0001) )  \state_ns_a2_0_0_a2_0_5[8]  (.A(
        pulse_meash_0_new_ready), .B(un1_i_cry_22_S), .C(
        un1_i_cry_23_S), .D(un1_i_cry_24_S), .Y(
        \state_ns_a2_0_0_a2_0_5[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_10 (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_9_net_1), .S(un1_i_cry_10_S), .Y(), .FCO(
        un1_i_cry_10_net_1));
    CFG4 #( .INIT(16'hBFFF) )  un38_clk_cry_30_RNILS9U_0 (.A(dir_net_1)
        , .B(FCCC_0_LOCK), .C(un38_clk_cry_30_net_1), .D(
        \state[2]_net_1 ), .Y(N_191_i_0_0));
    SLE \state[9]  (.D(\state[10]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[9]_net_1 ));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIMAN0K[5]  (.A(N_191_i_0), 
        .B(un46_clk_5), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[4] ), .S(\cr_angle_s[5] ), .Y(), .FCO(
        \cr_angle_cry[5] ));
    SLE en_timer (.D(\state[6]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_244_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(
        locator_control_0_en_timer));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_7 (.A(VCC_net_1), .B(
        un46_clk_7), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_6_net_1), .S(), .Y(), .FCO(un38_clk_cry_7_net_1));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_23 (.A(VCC_net_1), .B(
        un46_clk_23), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_22_net_1), .S(), .Y(), .FCO(un38_clk_cry_23_net_1)
        );
    CFG3 #( .INIT(8'h04) )  \state_RNO[2]  (.A(N_452_1), .B(
        \state[3]_net_1 ), .C(N_192), .Y(N_211_i_0));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_6 (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_5_net_1), .S(un1_i_cry_6_S), .Y(), .FCO(
        un1_i_cry_6_net_1));
    SLE \cr_angle[11]  (.D(\cr_angle_s[11] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_11));
    SLE \i[25]  (.D(\i_4_i_i_a3[25]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[25]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_1 (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_s_1_322_FCO), .S(un1_i_cry_1_S), .Y(), .FCO(
        un1_i_cry_1_net_1));
    CFG4 #( .INIT(16'hFFEC) )  \state_ns[8]  (.A(\state[3]_net_1 ), .B(
        \state[4]_net_1 ), .C(N_452_1), .D(N_192), .Y(
        \state_ns[8]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[10]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_10_S), .C(N_446), .D(N_481), .Y(N_242));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI3D6O91[20]  (.A(N_191_i_0)
        , .B(un46_clk_20), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[19] ), .S(\cr_angle_s[20] ), .Y(), .FCO(
        \cr_angle_cry[20] ));
    CFG4 #( .INIT(16'hFEFF) )  un1_state_8_0_0_a2_RNIMPV61 (.A(
        \state[9]_net_1 ), .B(\state[0]_net_1 ), .C(\state[3]_net_1 ), 
        .D(N_503), .Y(N_243_i_0));
    CFG4 #( .INIT(16'h4CCC) )  \state_RNO[6]  (.A(N_449_5), .B(
        \state[7]_net_1 ), .C(N_449_9), .D(un1_state_8_0_0_o2_net_1), 
        .Y(N_204_i_0));
    SLE \i[15]  (.D(N_462), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[15]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_26 (.A(VCC_net_1), .B(
        un46_clk_26), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_25_net_1), .S(), .Y(), .FCO(un38_clk_cry_26_net_1)
        );
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIS8BLM1[29]  (.A(N_191_i_0)
        , .B(un46_clk_29), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[28] ), .S(\cr_angle_s[29] ), .Y(), .FCO(
        \cr_angle_cry[29] ));
    ARI1 #( .INIT(20'h5AA55) )  un46_clk_cry_2 (.A(un46_clk_2), .B(
        \st_angle[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_1_net_1), .S(), .Y(), .FCO(un46_clk_cry_2_net_1));
    SLE \cr_angle[13]  (.D(\cr_angle_s[13] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_13));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_22 (.A(VCC_net_1), .B(
        un46_clk_22), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_21_net_1), .S(), .Y(), .FCO(un46_clk_cry_22_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[7]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_7_S), .C(N_446), .D(N_481), .Y(N_456));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_7 (.A(VCC_net_1), .B(
        un46_clk_7), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_6_net_1), .S(), .Y(), .FCO(un46_clk_cry_7_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_cr_angle_1_sqmuxa_0_0 (.A(over_net_1), 
        .B(\state[1]_net_1 ), .C(N_291), .Y(
        un1_cr_angle_1_sqmuxa_0_0_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNINJ0HI[4]  (.A(N_191_i_0), 
        .B(un46_clk_4), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[3] ), .S(\cr_angle_s[4] ), .Y(), .FCO(
        \cr_angle_cry[4] ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_5 (.A(VCC_net_1), .B(
        un46_clk_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_4_net_1), .S(), .Y(), .FCO(un38_clk_cry_5_net_1));
    ARI1 #( .INIT(20'h5CCAA) )  un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83 
        (.A(VCC_net_1), .B(N_191_i_0_0), .C(N_451_i_0), .D(GND_net_1), 
        .FCI(cr_angle_lcry_cy), .S(), .Y(
        un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y), .FCO(cr_angle));
    CFG4 #( .INIT(16'h5554) )  \i_4_i_i_a3[0]  (.A(\i[0]_net_1 ), .B(
        \state[3]_net_1 ), .C(N_446), .D(N_481), .Y(N_230));
    SLE \i[22]  (.D(\i_4_i_i_a3[22]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[22]_net_1 ));
    SLE \cr_angle[26]  (.D(\cr_angle_s[26] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_26));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_10 (.A(VCC_net_1), .B(
        un46_clk_10), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_9_net_1), .S(), .Y(), .FCO(un46_clk_cry_10_net_1));
    CFG4 #( .INIT(16'hC400) )  \state_ns_0_a3[11]  (.A(\i[21]_net_1 ), 
        .B(\state[0]_net_1 ), .C(N_491), .D(N_258), .Y(N_481));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI0T59U[12]  (.A(N_191_i_0), 
        .B(un46_clk_12), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[11] ), .S(\cr_angle_s[12] ), .Y(), .FCO(
        \cr_angle_cry[12] ));
    SLE \cr_angle[30]  (.D(\cr_angle_s[30] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_30));
    SLE \cr_angle[25]  (.D(\cr_angle_s[25] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_25));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_4 (.A(VCC_net_1), .B(
        un46_clk_4), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_3_net_1), .S(), .Y(), .FCO(un46_clk_cry_4_net_1));
    CFG4 #( .INIT(16'h7F77) )  \state_ns_i_0_0_o2_4[3]  (.A(
        \i[8]_net_1 ), .B(\i[7]_net_1 ), .C(\i[6]_net_1 ), .D(N_109), 
        .Y(N_116));
    CFG3 #( .INIT(8'h10) )  \state_ns_i_0_0_a2[3]  (.A(\i[20]_net_1 ), 
        .B(\i[19]_net_1 ), .C(N_120), .Y(N_491));
    CFG4 #( .INIT(16'hDFFF) )  un1_state_8_0_0_o2 (.A(\i[4]_net_1 ), 
        .B(un1_state_8_0_0_o2_2_net_1), .C(\i[6]_net_1 ), .D(
        \i[5]_net_1 ), .Y(un1_state_8_0_0_o2_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI01KBI1[26]  (.A(N_191_i_0)
        , .B(un46_clk_26), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[25] ), .S(\cr_angle_s[26] ), .Y(), .FCO(
        \cr_angle_cry[26] ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_28 (.A(VCC_net_1), .B(
        un46_clk_28), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_27_net_1), .S(), .Y(), .FCO(un38_clk_cry_28_net_1)
        );
    SLE \i[2]  (.D(N_232), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    SLE \i[12]  (.D(N_459), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_15 (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_14_net_1), .S(un1_i_cry_15_S), .Y(), .FCO(
        un1_i_cry_15_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNINI9A81[19]  (.A(N_191_i_0)
        , .B(un46_clk_19), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[18] ), .S(\cr_angle_s[19] ), .Y(), .FCO(
        \cr_angle_cry[19] ));
    SLE \state[8]  (.D(N_201_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[8]_net_1 ));
    CFG2 #( .INIT(4'h1) )  un1_state_8_0_0_a2 (.A(\state[8]_net_1 ), 
        .B(\state[7]_net_1 ), .Y(N_503));
    CFG2 #( .INIT(4'hE) )  en_timer_RNO (.A(\state[4]_net_1 ), .B(
        \state[6]_net_1 ), .Y(N_244_i_0));
    SLE \cr_angle[9]  (.D(\cr_angle_s[9] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_9));
    SLE \i[20]  (.D(N_467), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[20]_net_1 ));
    SLE \i[30]  (.D(\i_4_i_i_a3[30]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[30]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_14 (.A(VCC_net_1), .B(
        un46_clk_14), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_13_net_1), .S(), .Y(), .FCO(un46_clk_cry_14_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_9 (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_8_net_1), .S(un1_i_cry_9_S), .Y(), .FCO(
        un1_i_cry_9_net_1));
    SLE \state[3]  (.D(\state_ns[8]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[3]_net_1 ));
    SLE \fn_angle[2]  (.D(BT_module_0_data_buf[6]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un38_clk_2));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_18 (.A(VCC_net_1), .B(
        un46_clk_18), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_17_net_1), .S(), .Y(), .FCO(un46_clk_cry_18_net_1)
        );
    SLE over (.D(over_1_sqmuxa), .CLK(FCCC_0_GL0), .EN(
        un1_angle_0_sqmuxa_0_0_net_1), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(over_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_18 (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_17_net_1), .S(un1_i_cry_18_S), .Y(), .FCO(
        un1_i_cry_18_net_1));
    SLE \i[10]  (.D(N_242), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un1_state_8_0_0_a3_10_3 (.A(
        \i[20]_net_1 ), .B(\i[19]_net_1 ), .C(\i[12]_net_1 ), .D(
        \i[11]_net_1 ), .Y(un1_state_8_0_0_a3_10_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_14 (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_13_net_1), .S(un1_i_cry_14_S), .Y(), .FCO(
        un1_i_cry_14_net_1));
    SLE \i[6]  (.D(N_455), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_29 (.A(VCC_net_1), .B(
        un46_clk_29), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_28_net_1), .S(), .Y(), .FCO(un38_clk_cry_29_net_1)
        );
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_11 (.A(VCC_net_1), .B(
        un46_clk_11), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_10_net_1), .S(), .Y(), .FCO(un38_clk_cry_11_net_1)
        );
    SLE \i[29]  (.D(\i_4_i_i_a3[29]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[29]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \state_ns_0[4]  (.A(N_446), .B(
        \state[8]_net_1 ), .Y(\state_ns[4] ));
    SLE \fn_angle[3]  (.D(BT_module_0_data_buf[7]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un38_clk_3));
    SLE \st_angle[1]  (.D(BT_module_0_data_buf[1]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \st_angle[1]_net_1 ));
    SLE \i[4]  (.D(N_234), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_27 (.A(VCC_net_1), .B(
        un46_clk_27), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_26_net_1), .S(), .Y(), .FCO(un46_clk_cry_27_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_17 (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_16_net_1), .S(un31_clklto17), .Y(), .FCO(
        un1_i_cry_17_net_1));
    ARI1 #( .INIT(20'h4FDDD) )  un1_cr_angle_1_sqmuxa_0_0_a2_RNIN8VQ1 
        (.A(un38_clk_cry_30_net_1), .B(FCCC_0_LOCK), .C(N_229), .D(
        N_291), .FCI(VCC_net_1), .S(), .Y(), .FCO(cr_angle_lcry_cy));
    SLE \cr_angle[3]  (.D(\cr_angle_s[3] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_3));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_16 (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_15_net_1), .S(un1_i_cry_16_S), .Y(), .FCO(
        un1_i_cry_16_net_1));
    CFG4 #( .INIT(16'h5755) )  \state_ns_i_0_0_o2_2[3]  (.A(
        \i[13]_net_1 ), .B(\i[12]_net_1 ), .C(\i[11]_net_1 ), .D(N_117)
        , .Y(N_118));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIPLRFO[8]  (.A(N_191_i_0), 
        .B(un46_clk_8), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[7] ), .S(\cr_angle_s[8] ), .Y(), .FCO(
        \cr_angle_cry[8] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_22 (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_21_net_1), .S(un1_i_cry_22_S), .Y(), .FCO(
        un1_i_cry_22_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIUGL041[16]  (.A(N_191_i_0)
        , .B(un46_clk_16), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[15] ), .S(\cr_angle_s[16] ), .Y(), .FCO(
        \cr_angle_cry[16] ));
    SLE \i[19]  (.D(N_466), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[19]_net_1 ));
    SLE \cr_angle[17]  (.D(\cr_angle_s[17] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_17));
    SLE \st_angle[0]  (.D(BT_module_0_data_buf[0]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \st_angle[0]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[20]  (.A(\state[3]_net_1 ), 
        .B(un31_clklto20), .C(N_446), .D(N_481), .Y(N_467));
    SLE \cr_angle[12]  (.D(\cr_angle_s[12] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_12));
    SLE \cr_angle[19]  (.D(\cr_angle_s[19] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_19));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_10 (.A(VCC_net_1), .B(
        un46_clk_10), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_9_net_1), .S(), .Y(), .FCO(un38_clk_cry_10_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_20 (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_19_net_1), .S(un31_clklto20), .Y(), .FCO(
        un1_i_cry_20_net_1));
    CFG4 #( .INIT(16'h0080) )  \state_ns_a2_0_0_a3_0_7[8]  (.A(
        \state[3]_net_1 ), .B(\i[0]_net_1 ), .C(
        \state_ns_a2_0_0_a3_0_5[8]_net_1 ), .D(un31_clklto17), .Y(
        \state_ns_a2_0_0_a3_0_7[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_s_1_322 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(un1_i_s_1_322_FCO));
    SLE \angle1[0]  (.D(un46_clk_0), .CLK(FCCC_0_GL0), .EN(
        \state[4]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        locator_control_0_angle1[0]));
    CFG2 #( .INIT(4'hE) )  \state_ns_0[11]  (.A(N_481), .B(N_234_0), 
        .Y(\state_ns[11] ));
    SLE \i[24]  (.D(\i_4_i_i_a3[24]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[24]_net_1 ));
    SLE \cr_angle[5]  (.D(\cr_angle_s[5] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_5));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_2 (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_1_net_1), .S(un1_i_cry_2_S), .Y(), .FCO(
        un1_i_cry_2_net_1));
    CFG4 #( .INIT(16'h0001) )  un1_state_8_0_0_a3_10_2 (.A(
        \i[18]_net_1 ), .B(\i[13]_net_1 ), .C(\i[10]_net_1 ), .D(
        \i[9]_net_1 ), .Y(un1_state_8_0_0_a3_10_2_net_1));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_15 (.A(VCC_net_1), .B(
        un46_clk_15), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_14_net_1), .S(), .Y(), .FCO(un46_clk_cry_15_net_1)
        );
    SLE \cr_angle[24]  (.D(\cr_angle_s[24] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_24));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIM2EGL[6]  (.A(N_191_i_0), 
        .B(un46_clk_6), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[5] ), .S(\cr_angle_s[6] ), .Y(), .FCO(
        \cr_angle_cry[6] ));
    CFG3 #( .INIT(8'hF8) )  un1_angle_0_sqmuxa_0_0 (.A(over_net_1), .B(
        \state[1]_net_1 ), .C(over_1_sqmuxa), .Y(
        un1_angle_0_sqmuxa_0_0_net_1));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_20 (.A(VCC_net_1), .B(
        un46_clk_20), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_19_net_1), .S(), .Y(), .FCO(un46_clk_cry_20_net_1)
        );
    CFG4 #( .INIT(16'h1000) )  \state_ns_a2_0_a2[4]  (.A(\i[24]_net_1 )
        , .B(\i[26]_net_1 ), .C(\state_ns_a2_0_a2_5[4]_net_1 ), .D(
        \state_ns_a2_0_a2_4[4]_net_1 ), .Y(N_258));
    CFG3 #( .INIT(8'h01) )  \state_ns_a2_0_a2_2[4]  (.A(\i[16]_net_1 ), 
        .B(\i[15]_net_1 ), .C(\i[14]_net_1 ), .Y(N_59));
    SLE \i[14]  (.D(N_461), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    SLE \angle1[3]  (.D(un46_clk_3), .CLK(FCCC_0_GL0), .EN(
        \state[4]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        locator_control_0_angle1[3]));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_9 (.A(VCC_net_1), .B(
        un46_clk_9), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_8_net_1), .S(), .Y(), .FCO(un38_clk_cry_9_net_1));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[12]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_12_S), .C(N_446), .D(N_481), .Y(N_459));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[17]  (.A(\state[3]_net_1 ), 
        .B(un31_clklto17), .C(N_446), .D(N_481), .Y(N_464));
    SLE \fn_angle[0]  (.D(BT_module_0_data_buf[4]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un38_clk_0));
    SLE \state[2]  (.D(N_211_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[11]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_11_S), .C(N_446), .D(N_481), .Y(N_458));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_3 (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_2_net_1), .S(un1_i_cry_3_S), .Y(), .FCO(
        un1_i_cry_3_net_1));
    SLE en_sonar (.D(\state[8]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_state_8_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(TRIG_c));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_27 (.A(VCC_net_1), .B(
        un46_clk_27), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_26_net_1), .S(), .Y(), .FCO(un38_clk_cry_27_net_1)
        );
    SLE \state[1]  (.D(\state[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    SLE \cr_angle[28]  (.D(\cr_angle_s[28] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_28));
    CFG2 #( .INIT(4'h1) )  un1_state_8_0_0_a3_5 (.A(\i[21]_net_1 ), .B(
        \i[17]_net_1 ), .Y(N_449_5));
    SLE \i[5]  (.D(N_235), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    SLE \i[8]  (.D(N_457), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_24 (.A(VCC_net_1), .B(
        un46_clk_24), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_23_net_1), .S(), .Y(), .FCO(un46_clk_cry_24_net_1)
        );
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_19 (.A(VCC_net_1), .B(
        un46_clk_19), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_18_net_1), .S(), .Y(), .FCO(un46_clk_cry_19_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[6]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_6_S), .C(N_446), .D(N_481), .Y(N_455));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIGGHE51[17]  (.A(N_191_i_0)
        , .B(un46_clk_17), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[16] ), .S(\cr_angle_s[17] ), .Y(), .FCO(
        \cr_angle_cry[17] ));
    CFG4 #( .INIT(16'h08CC) )  \state_RNO[8]  (.A(\i[21]_net_1 ), .B(
        \state[0]_net_1 ), .C(N_491), .D(N_258), .Y(N_201_i_0));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_22 (.A(VCC_net_1), .B(
        un46_clk_22), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_21_net_1), .S(), .Y(), .FCO(un38_clk_cry_22_net_1)
        );
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_28 (.A(VCC_net_1), .B(
        un46_clk_28), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_27_net_1), .S(), .Y(), .FCO(un46_clk_cry_28_net_1)
        );
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_8 (.A(VCC_net_1), .B(
        un46_clk_8), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_7_net_1), .S(), .Y(), .FCO(un38_clk_cry_8_net_1));
    SLE \cr_angle[7]  (.D(\cr_angle_s[7] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_7));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_25 (.A(VCC_net_1), .B(
        \i[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_24_net_1), .S(un1_i_cry_25_S), .Y(), .FCO(
        un1_i_cry_25_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un38_clk_cry_1 (.A(un38_clk_1), .B(
        un46_clk_1), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_0_net_1), .S(), .Y(), .FCO(un38_clk_cry_1_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNID2T1E1[23]  (.A(N_191_i_0)
        , .B(un46_clk_23), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[22] ), .S(\cr_angle_s[23] ), .Y(), .FCO(
        \cr_angle_cry[23] ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_16 (.A(VCC_net_1), .B(
        un46_clk_16), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_15_net_1), .S(), .Y(), .FCO(un46_clk_cry_16_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[16]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_16_S), .C(N_446), .D(N_481), .Y(N_463));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[9]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_9_S), .C(N_446), .D(N_481), .Y(N_241));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIJ2HPJ1[27]  (.A(N_191_i_0)
        , .B(un46_clk_27), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[26] ), .S(\cr_angle_s[27] ), .Y(), .FCO(
        \cr_angle_cry[27] ));
    SLE \st_angle[3]  (.D(BT_module_0_data_buf[3]), .CLK(FCCC_0_GL0), 
        .EN(fn_angle_0_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \st_angle[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_13 (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_12_net_1), .S(un1_i_cry_13_S), .Y(), .FCO(
        un1_i_cry_13_net_1));
    SLE \state[11]  (.D(N_195_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[11]_net_1 ));
    CFG4 #( .INIT(16'h777F) )  un1_state_8_0_0_o2_2 (.A(\i[8]_net_1 ), 
        .B(\i[7]_net_1 ), .C(\i[3]_net_1 ), .D(\i[2]_net_1 ), .Y(
        un1_state_8_0_0_o2_2_net_1));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_6 (.A(VCC_net_1), .B(
        un46_clk_6), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_5_net_1), .S(), .Y(), .FCO(un38_clk_cry_6_net_1));
    SLE \i[3]  (.D(N_233), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_28 (.A(VCC_net_1), .B(
        \i[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_27_net_1), .S(un1_i_cry_28_S), .Y(), .FCO(
        un1_i_cry_28_net_1));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIJ2ARS[11]  (.A(N_191_i_0), 
        .B(un46_clk_11), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[10] ), .S(\cr_angle_s[11] ), .Y(), .FCO(
        \cr_angle_cry[11] ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_5 (.A(VCC_net_1), .B(
        un46_clk_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_4_net_1), .S(), .Y(), .FCO(un46_clk_cry_5_net_1));
    CFG4 #( .INIT(16'h7500) )  \state_ns_i_0_0_a3[9]  (.A(
        un31_clklto21), .B(un31_clklto20), .C(N_114), .D(N_311), .Y(
        N_452_1));
    CFG4 #( .INIT(16'h8000) )  \state_ns_a2_0_0_a3_0[8]  (.A(
        \state_ns_a2_0_0_a3_0_7[8]_net_1 ), .B(N_311), .C(N_316), .D(
        \state_ns_a2_0_0_a3_0_6[8]_net_1 ), .Y(N_192));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNINR40N[7]  (.A(N_191_i_0), 
        .B(un46_clk_7), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), .FCI(
        \cr_angle_cry[6] ), .S(\cr_angle_s[7] ), .Y(), .FCO(
        \cr_angle_cry[7] ));
    SLE \cr_angle[4]  (.D(\cr_angle_s[4] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_4));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_24 (.A(VCC_net_1), .B(
        \i[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_23_net_1), .S(un1_i_cry_24_S), .Y(), .FCO(
        un1_i_cry_24_net_1));
    ARI1 #( .INIT(20'h51BE4) )  \st_angle_RNIB8ELC[2]  (.A(N_191_i_0), 
        .B(un1_cr_angle_1_sqmuxa_0_0_a2_RNI1LN83_Y), .C(
        \st_angle[2]_net_1 ), .D(un46_clk_2), .FCI(\cr_angle_cry[1] ), 
        .S(\cr_angle_s[2] ), .Y(), .FCO(\cr_angle_cry[2] ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_25 (.A(VCC_net_1), .B(
        un46_clk_25), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_24_net_1), .S(), .Y(), .FCO(un38_clk_cry_25_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_11 (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_10_net_1), .S(un1_i_cry_11_S), .Y(), .FCO(
        un1_i_cry_11_net_1));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_14 (.A(VCC_net_1), .B(
        un46_clk_14), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_13_net_1), .S(), .Y(), .FCO(un38_clk_cry_14_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_27 (.A(VCC_net_1), .B(
        \i[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_26_net_1), .S(un1_i_cry_27_S), .Y(), .FCO(
        un1_i_cry_27_net_1));
    CFG4 #( .INIT(16'hB8F0) )  \st_angle_RNI7D8K[0]  (.A(
        \st_angle[0]_net_1 ), .B(FCCC_0_LOCK), .C(un46_clk_0), .D(
        \state[10]_net_1 ), .Y(\cr_angle_lxu;_0[0] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_26 (.A(VCC_net_1), .B(
        \i[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_25_net_1), .S(un1_i_cry_26_S), .Y(), .FCO(
        un1_i_cry_26_net_1));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[13]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_13_S), .C(N_446), .D(N_481), .Y(N_460));
    SLE \i[1]  (.D(N_231), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[3]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_3_S), .C(N_446), .D(N_481), .Y(N_233));
    SLE \cr_angle[0]  (.D(\cr_angle_s[0] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_0));
    SLE \cr_angle[20]  (.D(\cr_angle_s[20] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_20));
    SLE \i[28]  (.D(\i_4_i_i_a3[28]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[28]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_13 (.A(VCC_net_1), .B(
        un46_clk_13), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_12_net_1), .S(), .Y(), .FCO(un38_clk_cry_13_net_1)
        );
    CFG4 #( .INIT(16'h5DFF) )  \state_ns_a2_0_0_o2_0[8]  (.A(
        un1_i_cry_19_S), .B(N_112), .C(un31_clklto17), .D(
        un1_i_cry_18_S), .Y(N_114));
    CFG2 #( .INIT(4'h6) )  \cr_angle_qxu[0]  (.A(N_191_i_0), .B(
        \cr_angle_lxu;[0] ), .Y(\cr_angle_qxu[0]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  \state_ns_a2_0_0_a2_0[8]  (.A(
        un1_i_cry_29_S), .B(un1_i_s_30_S), .C(
        \state_ns_a2_0_0_a2_0_5[8]_net_1 ), .D(
        \state_ns_a2_0_0_a2_0_6[8]_net_1 ), .Y(N_311));
    SLE \cr_angle[16]  (.D(\cr_angle_s[16] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_16));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_25 (.A(VCC_net_1), .B(
        un46_clk_25), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_24_net_1), .S(), .Y(), .FCO(un46_clk_cry_25_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[4]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_4_S), .C(N_446), .D(N_481), .Y(N_234));
    SLE \cr_angle[15]  (.D(\cr_angle_s[15] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_15));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_19 (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_18_net_1), .S(un1_i_cry_19_S), .Y(), .FCO(
        un1_i_cry_19_net_1));
    CFG3 #( .INIT(8'h13) )  \state_ns_a2_0_0_a2_13[8]  (.A(
        un1_i_cry_7_S), .B(un31_clklto8), .C(un1_i_cry_6_S), .Y(N_482));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[22]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_22_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[22]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[27]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_27_S), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[27]_net_1 ));
    SLE \i[18]  (.D(N_465), .CLK(FCCC_0_GL0), .EN(N_243_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[18]_net_1 ));
    SLE \cr_angle[1]  (.D(\cr_angle_s[1] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(un46_clk_1));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[21]  (.A(\state[3]_net_1 ), 
        .B(un31_clklto21), .C(N_446), .D(N_481), .Y(
        \i_4_i_i_a3[21]_net_1 ));
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[14]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_14_S), .C(N_446), .D(N_481), .Y(N_461));
    ARI1 #( .INIT(20'h45500) )  un38_clk_cry_16 (.A(VCC_net_1), .B(
        un46_clk_16), .C(GND_net_1), .D(GND_net_1), .FCI(
        un38_clk_cry_15_net_1), .S(), .Y(), .FCO(un38_clk_cry_16_net_1)
        );
    CFG4 #( .INIT(16'hCCC8) )  \i_4_i_i_a3[19]  (.A(\state[3]_net_1 ), 
        .B(un1_i_cry_19_S), .C(N_446), .D(N_481), .Y(N_466));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNI3HDS61[18]  (.A(N_191_i_0)
        , .B(un46_clk_18), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[17] ), .S(\cr_angle_s[18] ), .Y(), .FCO(
        \cr_angle_cry[18] ));
    ARI1 #( .INIT(20'h65500) )  un46_clk_cry_13 (.A(VCC_net_1), .B(
        un46_clk_13), .C(GND_net_1), .D(GND_net_1), .FCI(
        un46_clk_cry_12_net_1), .S(), .Y(), .FCO(un46_clk_cry_13_net_1)
        );
    CFG3 #( .INIT(8'h08) )  un1_angle_0_sqmuxa_0_0_a3_0 (.A(dir_net_1), 
        .B(\state[2]_net_1 ), .C(un46_clk_cry_30_net_1), .Y(
        over_1_sqmuxa));
    ARI1 #( .INIT(20'h5D52A) )  \cr_angle_RNIT0QFF1[24]  (.A(N_191_i_0)
        , .B(un46_clk_24), .C(FCCC_0_LOCK), .D(\state[10]_net_1 ), 
        .FCI(\cr_angle_cry[23] ), .S(\cr_angle_s[24] ), .Y(), .FCO(
        \cr_angle_cry[24] ));
    SLE \i[26]  (.D(\i_4_i_i_a3[26]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_243_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\i[26]_net_1 ));
    
endmodule


module time_sender(
       locator_control_0_angle1,
       pulse_meash_0_tim,
       time_sender_0_data_out_0,
       time_sender_0_data_out_1,
       time_sender_0_data_out_2,
       time_sender_0_data_out_3,
       time_sender_0_data_out_5,
       LED_3_c,
       LED_3_c_i_0,
       FCCC_0_GL0,
       FCCC_0_LOCK,
       pulse_meash_0_new_ready,
       COREUART_0_TXRDY
    );
input  [3:0] locator_control_0_angle1;
input  [13:0] pulse_meash_0_tim;
output time_sender_0_data_out_0;
output time_sender_0_data_out_1;
output time_sender_0_data_out_2;
output time_sender_0_data_out_3;
output time_sender_0_data_out_5;
output LED_3_c;
output LED_3_c_i_0;
input  FCCC_0_GL0;
input  FCCC_0_LOCK;
input  pulse_meash_0_new_ready;
input  COREUART_0_TXRDY;

    wire \valu[6]_net_1 , VCC_net_1, \un1_time1[6]_net_1 , 
        un1_rst_n_inv_i_a3_net_1, GND_net_1, \valu[7]_net_1 , 
        \un1_time1[7]_net_1 , \valu[8]_net_1 , \un1_time1[8]_net_1 , 
        \valu[9]_net_1 , \un1_time1[9]_net_1 , \valu[10]_net_1 , 
        \un1_time1[10]_net_1 , \valu[11]_net_1 , \valu_RNO[11]_net_1 , 
        \valu[12]_net_1 , \valu_RNO[12]_net_1 , \valu[13]_net_1 , 
        \un1_time1[13]_net_1 , \data_out_1[0] , data_out_0_sqmuxa, 
        \data_out_1[1] , \data_out_1[2] , \data_out_1[3] , 
        \data_out_1[5] , \valu[0]_net_1 , \un1_time1[0]_net_1 , 
        \valu[1]_net_1 , \un1_time1[1]_net_1 , \valu[2]_net_1 , 
        \un1_time1[2]_net_1 , \valu[3]_net_1 , \un1_time1[3]_net_1 , 
        \valu[4]_net_1 , \un1_time1[4]_net_1 , \valu[5]_net_1 , 
        \un1_time1[5]_net_1 , \k[0]_net_1 , N_87_i_0, \k[1]_net_1 , 
        \un24_k_v[0]_net_1 , \k[2]_net_1 , \un24_k_v[1]_net_1 , 
        \k[3]_net_1 , \SUM[3] , \k[5] , \buff_1[0]_net_1 , 
        \un1_angle[0]_net_1 , un1_rst_n_inv_2_i_0_net_1, 
        \buff_1[1]_net_1 , \un1_angle[1]_net_1 , \buff_1[2]_net_1 , 
        \un1_angle[2]_net_1 , \buff_1[3]_net_1 , \un1_angle[3]_net_1 , 
        \buff_1[5] , \un1_angle[4]_net_1 , \buff_3[1]_net_1 , 
        buff_3_1_sqmuxa_net_1, \buff_3[2]_net_1 , \buff_3[3]_net_1 , 
        \buff_3[5] , \buff_2[0]_net_1 , buff_2_1_sqmuxa_1_net_1, 
        \buff_2[1]_net_1 , \buff_2[2]_net_1 , \buff_2[3]_net_1 , 
        \buff_2[5] , \buff_5[2]_net_1 , buff_5_1_sqmuxa_net_1, 
        \buff_5[3]_net_1 , \buff_5[5] , \buff_4[0]_net_1 , 
        buff_4_1_sqmuxa_net_1, \buff_4[1]_net_1 , \buff_4[2]_net_1 , 
        \buff_4[3]_net_1 , \buff_4[5] , \buff_3[0]_net_1 , 
        \buff_5[0]_net_1 , \buff_5[1]_net_1 , \buff_0[5] , 
        buff_0_1_sqmuxa, N_139_i_0, N_445_i_0, \buff_0[0]_net_1 , 
        \buff_0[1]_net_1 , \buff_0[2]_net_1 , \buff_0[3]_net_1 , 
        \state[6]_net_1 , \state_ns[0] , \state[5]_net_1 , N_85_i_0, 
        \state[4]_net_1 , \state[3]_net_1 , N_10_i_0, \state[2]_net_1 , 
        N_431_i_0, \state[1]_net_1 , N_84_tz_i, \state[0]_net_1 , 
        \state_ns[6] , \i[0]_net_1 , \i_lm[0] , N_84_i_0, \i[1]_net_1 , 
        \i_lm[1] , \i[2]_net_1 , \i_lm[2] , \i[3]_net_1 , \i_lm[3] , 
        \i[4]_net_1 , \i_lm[4] , \i[5]_net_1 , \i_lm[5] , \i[6]_net_1 , 
        \i_lm[6] , \i[7]_net_1 , \i_lm[7] , \i[8]_net_1 , \i_lm[8] , 
        \i[9]_net_1 , \i_lm[9] , \i[10]_net_1 , \i_lm[10] , 
        \i[11]_net_1 , \i_lm[11] , \i[12]_net_1 , \i_lm[12] , 
        \i[13]_net_1 , \i_lm[13] , \i[14]_net_1 , \i_lm[14] , 
        \i[15]_net_1 , \i_lm[15] , \i[16]_net_1 , \i_lm[16] , 
        \i[17]_net_1 , \i_lm[17] , \i[18]_net_1 , \i_lm[18] , 
        \i[19]_net_1 , \i_lm[19] , \i[20]_net_1 , \i_lm[20] , 
        \i[21]_net_1 , \i_lm[21] , \i[22]_net_1 , \i_lm[22] , 
        \i[23]_net_1 , \i_lm[23] , \i[24]_net_1 , \i_lm[24] , 
        \i[25]_net_1 , \i_lm[25] , \i_cry[0]_net_1 , \i_cry_Y_0[0] , 
        \i_cry[1]_net_1 , \i_s[1] , \i_cry[2]_net_1 , \i_s[2] , 
        \i_cry[3]_net_1 , \i_s[3] , \i_cry[4]_net_1 , \i_s[4] , 
        \i_cry[5]_net_1 , \i_s[5] , \i_cry[6]_net_1 , \i_s[6] , 
        \i_cry[7]_net_1 , \i_s[7] , \i_cry[8]_net_1 , \i_s[8] , 
        \i_cry[9]_net_1 , \i_s[9] , \i_cry[10]_net_1 , \i_s[10] , 
        \i_cry[11]_net_1 , \i_s[11] , \i_cry[12]_net_1 , \i_s[12] , 
        \i_cry[13]_net_1 , \i_s[13] , \i_cry[14]_net_1 , \i_s[14] , 
        \i_cry[15]_net_1 , \i_s[15] , \i_cry[16]_net_1 , \i_s[16] , 
        \i_cry[17]_net_1 , \i_s[17] , \i_cry[18]_net_1 , \i_s[18] , 
        \i_cry[19]_net_1 , \i_s[19] , \i_cry[20]_net_1 , \i_s[20] , 
        \i_cry[21]_net_1 , \i_s[21] , \i_cry[22]_net_1 , \i_s[22] , 
        \i_cry[23]_net_1 , \i_s[23] , \i_s[25]_net_1 , 
        \i_cry[24]_net_1 , \i_s[24] , un1_i_s_1_323_FCO, 
        un1_i_cry_1_net_1, un15_clklto1, un1_i_cry_2_net_1, 
        un15_clklto2, un1_i_cry_3_net_1, un1_i_cry_3_S_0, 
        un1_i_cry_4_net_1, un1_i_cry_4_S_0, un1_i_cry_5_net_1, 
        un1_i_cry_5_S_0, un1_i_cry_6_net_1, un1_i_cry_6_S_0, 
        un1_i_cry_7_net_1, un1_i_cry_7_S_0, un1_i_cry_8_net_1, 
        un1_i_cry_8_S, un1_i_cry_9_net_1, un1_i_cry_9_S_0, 
        un1_i_cry_10_net_1, un1_i_cry_10_S_0, un1_i_cry_11_net_1, 
        un1_i_cry_11_S_0, un1_i_cry_12_net_1, un1_i_cry_12_S_0, 
        un1_i_cry_13_net_1, un1_i_cry_13_S_0, un1_i_cry_14_net_1, 
        un1_i_cry_14_S_0, un1_i_cry_15_net_1, un1_i_cry_15_S_0, 
        un1_i_cry_16_net_1, un1_i_cry_16_S_0, un1_i_cry_17_net_1, 
        un1_i_cry_17_S, un1_i_cry_18_net_1, un1_i_cry_18_S_0, 
        un1_i_cry_19_net_1, un1_i_cry_19_S_0, un1_i_cry_20_net_1, 
        un1_i_cry_20_S, un1_i_cry_21_net_1, un1_i_cry_21_S, 
        un1_i_cry_22_net_1, un1_i_cry_22_S_0, un1_i_cry_23_net_1, 
        un1_i_cry_23_S_0, un1_i_cry_24_net_1, un1_i_cry_24_S_0, 
        un1_i_cry_25_net_1, un1_i_cry_25_S_0, 
        \mult1_un215_sum_1_SUM[4] , mult1_un222_sum_1_CO1, 
        \mult1_un215_sum_1_SUM[1] , \mult1_un215_sum_1_SUM[2] , 
        mult1_un222_sum_1_CO3, \un1_clk_inv_i_0_o3[0]_net_1 , 
        un1_N_3_mux, \valu_RNICB5V[13]_net_1 , N_91, 
        \state_ns_i_a2[3]_net_1 , N_96, \mult1_un166_sum_1_SUM[2] , 
        mult1_un166_sum_1_CO3, un1_N_13_mux, un1_i4_mux, N_3560_i, 
        \mult1_un194_sum_1_SUM[2] , un1_m7_i_0_1, un1_N_8, un1_m7_i_0, 
        mult1_un201_sum_1_CO2_0_tz, mult1_un201_sum_1_ANC2, 
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42, un1_m9_1, 
        mult1_un187_sum_1_CO3_1_RNIDREF, \mult1_un194_sum_1_SUM_1[4] , 
        mult1_un194_sum_1_CO3_0_tz, \mult1_un187_sum_1_SUM[2] , 
        d_m2_3_0, \mult1_un187_sum_1_SUM[1] , 
        mult1_un194_sum_1_ANC3_0_1_1, \mult1_un187_sum_1_SUM[4] , 
        mult1_un194_sum_1_ANC3_0_1, mult1_un194_sum_1_CO3_0_tz_0_1, 
        mult1_un194_sum_1_CO3_0_tz_0_RNO, \mult1_un180_sum_1_SUM[1] , 
        mult1_un194_sum_1_CO3_0_tz_0_1_RNO, \mult1_un180_sum_1_SUM[4] , 
        \mult1_un180_sum_1_SUM[2] , un1_m8_1_1, 
        \mult1_un159_sum_1_SUM[4] , \mult1_un159_sum_1_SUM[1] , 
        \mult1_un159_sum_1_SUM[2] , un1_m8_1, 
        \data_out_1_5_am_1_1[4]_net_1 , \data_out_1_5_am[4]_net_1 , 
        \data_out_1_5_am_1_1[3]_net_1 , \data_out_1_5_am[3]_net_1 , 
        \data_out_1_5_am_1_1[2]_net_1 , \data_out_1_5_am[2]_net_1 , 
        \data_out_1_5_am_1_1[1]_net_1 , \data_out_1_5_am[1]_net_1 , 
        \data_out_1_5_am_1_1[0]_net_1 , \data_out_1_5_am[0]_net_1 , 
        \valu_RNINMIF[13]_net_1 , \valu_RNI32OE1[13]_net_1 , 
        \mult1_un159_sum_1_SUM_2_1[4] , \data_out_1_5_bm[4]_net_1 , 
        \data_out_1_5_bm[3]_net_1 , \data_out_1_5_bm[2]_net_1 , 
        \data_out_1_5_bm[1]_net_1 , \data_out_1_5_bm[0]_net_1 , 
        \valu_RNILKIF_0[11]_net_1 , \mult1_un201_sum_1_SUM_1[1] , 
        un1_N_5_i_2, mult1_un194_sum_1_CO2, 
        \mult1_un201_sum_1_SUM_2[4] , \mult1_un173_sum_1_SUM[2] , 
        \mult1_un166_sum_1_SUM_RNIQ5884[1] , mult1_un180_sum_1_CO3_1, 
        d_m12_0_a3_0, d_N_4_1, N_89, N_90, buff_2_1_sqmuxa_net_1, 
        \state_ns_i_a2_17[3]_net_1 , \state_ns_i_a2_16[3]_net_1 , 
        \state_ns_i_a2_15[3]_net_1 , \state_ns_i_a2_14[3]_net_1 , 
        \state_ns_i_a2_13[3]_net_1 , \state_ns_i_a2_12[3]_net_1 , 
        \state_ns_i_0_a2_16[5]_net_1 , \state_ns_i_0_a2_15[5]_net_1 , 
        \state_ns_i_0_a2_14[5]_net_1 , \state_ns_i_0_a2_13[5]_net_1 , 
        \state_ns_i_0_a2_12[5]_net_1 , \state_ns_0_a3_3[0]_net_1 , 
        \state_ns_i_0_a2_17[5]_net_1 , N_104, 
        \state_ns_i_a2_21[3]_net_1 , \state_ns_i_0_a2_21[5]_net_1 , 
        \state_ns_i_0_a2_20[5]_net_1 , N_93, N_144, N_95, un1_m5_i_0, 
        mult1_un159_sum_1_CO3, mult1_un159_sum_1_CO3_1_RNI1HJB3, 
        un1_N_5_i_1, \mult1_un166_sum_1_SUM[1] , un1_N_5_1, 
        \mult1_un159_sum_1_SUM_RNIM44K4[4] , mult1_un173_sum_1_CO1_0, 
        \mult1_un166_sum_1_SUM[4] , \mult1_un173_sum_1_SUM[1] , 
        mult1_un180_sum_1_CO3_2_0, un1_m2_5_0, un1_i3_mux_0_0_i, 
        mult1_un180_sum_1_CO3_a4, \mult1_un180_sum_1_SUM_0[3] , 
        mult1_un180_sum_1_CO3_0_0, mult1_un173_sum_1_CO2, 
        \mult1_un180_sum_1_SUM_2[4] , un1_i1_mux, 
        mult1_un180_sum_1_CO2, mult1_un187_sum_1_CO3_1_RNO, 
        \mult1_un187_sum_1_SUM_0[4] , mult1_un187_sum_1_CO2, 
        un1_m4_1_1, mult1_un187_sum_1_CO3_0, d_N_12_0, d_m1_2_0, 
        d_i5_mux, d_N_2_0, un1_N_7_0, un1_m8_i_0, 
        \mult1_un194_sum_1_SUM[1] , d_N_10, d_N_19, d_N_11_mux_0, 
        un1_N_7_mux_0, d_N_11_mux, d_N_13_mux, 
        mult1_un201_sum_1_CO3_0_tz_s_0_RNO, 
        mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK, d_N_20, un1_i6_mux, 
        mult1_un201_sum_1_CO2_0_d_0_RNO_0, 
        mult1_un201_sum_1_ANC3_0_RNO_0, un1_N_10_mux, d_i6_mux_1, 
        mult1_un215_sum_1_CO3_0_RNO_3, mult1_un201_sum_1_CO2_0_d, 
        mult1_un201_sum_1_ANC3, mult1_un201_sum_1_CO3_0_tz_s_0, 
        mult1_un201_sum_1_CO1, mult1_un201_sum_1_CO3_0_d, 
        \mult1_un201_sum_1_SUM[2] , mult1_un201_sum_1_CO3_0_c, 
        mult1_un201_sum_1_CO3_0_0_1, un1_i3_mux_0, 
        mult1_un201_sum_1_CO3, \mult1_un201_sum_1_SUM[4] , 
        mult1_un201_sum_1_CO3_0_c_RNI45FP3, un1_N_5_mux, 
        \mult1_un215_sum_1_SUM_0_0[4] , un1_m6_1_0, un1_m7_3_0, 
        \mult1_un208_sum_1_SUM[1] , un1_N_7_i, mult1_un208_sum_1_CO2, 
        un1_i5_mux_0, un1_i2_mux, mult1_un215_sum_1_ANC3_0_RNO_0, 
        mult1_un215_sum_1_CO3_0_RNO, \mult1_un215_sum_1_SUM_0[3] , 
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] , mult1_un215_sum_1_ANC3, 
        \mult1_un215_sum_1_SUM_1[3] , \mult1_un215_sum_1_SUM_0[4] , 
        mult1_un215_sum_1_CO3_0, mult1_un215_sum_1_CO3, 
        mult1_un215_sum_1_CO1, \un24_k_v_1[1]_net_1 , \SUM_1[3] , 
        mult1_un215_sum_1_CO2, \mult1_un215_sum_1_SUM[3] , 
        \mult1_un222_sum_1_SUM_0[4] , ANC2_m3, CO2;
    
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_0_a2_13[5]  (.A(
        \i[18]_net_1 ), .B(\i[9]_net_1 ), .C(\i[8]_net_1 ), .D(
        \i[5]_net_1 ), .Y(\state_ns_i_0_a2_13[5]_net_1 ));
    CFG2 #( .INIT(4'h9) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0_RNO  (
        .A(mult1_un194_sum_1_CO3_0_tz), .B(
        \mult1_un194_sum_1_SUM_1[4] ), .Y(
        mult1_un201_sum_1_CO3_0_tz_s_0_RNO));
    SLE \state[0]  (.D(\state_ns[6] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    CFG4 #( .INIT(16'h0026) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0_RNO_3  
        (.A(\valu[6]_net_1 ), .B(\mult1_un187_sum_1_SUM[1] ), .C(
        \mult1_un187_sum_1_SUM[2] ), .D(\mult1_un187_sum_1_SUM[4] ), 
        .Y(un1_i6_mux));
    SLE \valu[10]  (.D(\un1_time1[10]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[10]_net_1 ));
    CFG4 #( .INIT(16'hC6CC) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_SUM[4]  (.A(
        mult1_un180_sum_1_CO3_1), .B(\mult1_un180_sum_1_SUM_2[4] ), .C(
        mult1_un180_sum_1_CO3_a4), .D(mult1_un180_sum_1_CO3_0_0), .Y(
        \mult1_un180_sum_1_SUM[4] ));
    CFG2 #( .INIT(4'h9) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM[1]  (.A(
        \mult1_un187_sum_1_SUM[4] ), .B(d_N_4_1), .Y(
        \mult1_un194_sum_1_SUM[1] ));
    SLE \i[7]  (.D(\i_lm[7] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    CFG3 #( .INIT(8'h31) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_ANC3_0_1_1  (.A(
        \valu[5]_net_1 ), .B(\mult1_un187_sum_1_SUM[1] ), .C(
        \valu[6]_net_1 ), .Y(mult1_un194_sum_1_ANC3_0_1_1));
    SLE \i[16]  (.D(\i_lm[16] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[16]_net_1 ));
    CFG4 #( .INIT(16'hC0AF) )  \data_out_1_5_am[0]  (.A(
        \buff_5[0]_net_1 ), .B(\buff_4[0]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\data_out_1_5_am_1_1[0]_net_1 ), .Y(
        \data_out_1_5_am[0]_net_1 ));
    CFG2 #( .INIT(4'hE) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3  (.A(
        mult1_un215_sum_1_CO3_0), .B(mult1_un215_sum_1_ANC3), .Y(
        mult1_un215_sum_1_CO3));
    CFG4 #( .INIT(16'h2000) )  buff_5_1_sqmuxa (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(buff_2_1_sqmuxa_net_1), .D(\i[0]_net_1 ), .Y(
        buff_5_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'h9669) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM[1]  (.A(
        \valu[3]_net_1 ), .B(\valu[2]_net_1 ), .C(un1_i2_mux), .D(
        un1_m6_1_0), .Y(\mult1_un215_sum_1_SUM[1] ));
    CFG4 #( .INIT(16'hF0E4) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0  (.A(
        un1_N_7_i), .B(\valu[2]_net_1 ), .C(
        mult1_un215_sum_1_ANC3_0_RNO_0), .D(un1_m7_i_0), .Y(
        mult1_un215_sum_1_ANC3));
    CFG4 #( .INIT(16'h0004) )  \state_ns_i_0_a2_20[5]  (.A(
        \i[0]_net_1 ), .B(\state_ns_i_0_a2_17[5]_net_1 ), .C(
        \i[1]_net_1 ), .D(\i[2]_net_1 ), .Y(
        \state_ns_i_0_a2_20[5]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  un1_rst_n_inv_2_i_a3_0 (.A(\i[2]_net_1 )
        , .B(\i[1]_net_1 ), .C(buff_2_1_sqmuxa_net_1), .D(\i[0]_net_1 )
        , .Y(N_104));
    SLE \buff_0[3]  (.D(\k[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_0_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_0[3]_net_1 ));
    CFG3 #( .INIT(8'h2E) )  \un1_time1[5]  (.A(pulse_meash_0_tim[5]), 
        .B(\state[4]_net_1 ), .C(\mult1_un187_sum_1_SUM[4] ), .Y(
        \un1_time1[5]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[14]  (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[13]_net_1 ), .S(\i_s[14] ), .Y(), .FCO(
        \i_cry[14]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  \state_ns_i_0_a2_17[5]  (.A(
        \i[21]_net_1 ), .B(\state_ns_i_0_a2_12[5]_net_1 ), .C(
        \i[25]_net_1 ), .D(\i[24]_net_1 ), .Y(
        \state_ns_i_0_a2_17[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[24]  (.A(\i_s[24] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[24] ));
    SLE \i[21]  (.D(\i_lm[21] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[21]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM_1[1]  (.A(
        \mult1_un194_sum_1_SUM_1[4] ), .B(\mult1_un187_sum_1_SUM[4] ), 
        .C(\valu[4]_net_1 ), .D(\valu[5]_net_1 ), .Y(
        \mult1_un201_sum_1_SUM_1[1] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[20]  (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[19]_net_1 ), .S(\i_s[20] ), .Y(), .FCO(
        \i_cry[20]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_14[3]  (.A(
        un1_i_cry_11_S_0), .B(un1_i_cry_12_S_0), .C(un1_i_cry_13_S_0), 
        .D(un1_i_cry_14_S_0), .Y(\state_ns_i_a2_14[3]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \un1_angle[2]  (.A(
        locator_control_0_angle1[2]), .B(\k[2]_net_1 ), .C(
        \state[4]_net_1 ), .Y(\un1_angle[2]_net_1 ));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM[2]  (.A(
        mult1_un201_sum_1_CO1), .B(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .C(
        \mult1_un194_sum_1_SUM[1] ), .Y(\mult1_un201_sum_1_SUM[2] ));
    CFG4 #( .INIT(16'hF702) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO_3  (.A(
        \mult1_un187_sum_1_SUM[2] ), .B(d_N_2_0), .C(d_N_12_0), .D(
        \mult1_un194_sum_1_SUM_1[4] ), .Y(d_N_13_mux));
    SLE \buff_4[1]  (.D(\k[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_4_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_4[1]_net_1 ));
    SLE \k[1]  (.D(\un24_k_v[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_87_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\k[1]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_ns[0]  (.A(
        \data_out_1_5_am[0]_net_1 ), .B(\i[1]_net_1 ), .C(
        \data_out_1_5_bm[0]_net_1 ), .Y(\data_out_1[0] ));
    SLE \i[0]  (.D(\i_lm[0] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \state_ns_i_0_a2_21[5]  (.A(
        \state_ns_i_0_a2_16[5]_net_1 ), .B(
        \state_ns_i_0_a2_15[5]_net_1 ), .C(
        \state_ns_i_0_a2_14[5]_net_1 ), .D(
        \state_ns_i_0_a2_13[5]_net_1 ), .Y(
        \state_ns_i_0_a2_21[5]_net_1 ));
    SLE \i[11]  (.D(\i_lm[11] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    CFG4 #( .INIT(16'h4644) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM_RNITTTU[2]  (.A(
        \mult1_un166_sum_1_SUM[2] ), .B(mult1_un166_sum_1_CO3), .C(
        \valu[9]_net_1 ), .D(\valu[8]_net_1 ), .Y(un1_i4_mux));
    CFG4 #( .INIT(16'h0001) )  \state_ns_0_a3_3[0]  (.A(
        \state[1]_net_1 ), .B(\state[5]_net_1 ), .C(\state[3]_net_1 ), 
        .D(\state[2]_net_1 ), .Y(\state_ns_0_a3_3[0]_net_1 ));
    SLE \state[6]  (.D(\state_ns[0] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[6]_net_1 ));
    CFG4 #( .INIT(16'hAE00) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_CO3_1  (.A(
        \mult1_un180_sum_1_SUM[2] ), .B(\mult1_un180_sum_1_SUM[1] ), 
        .C(un1_i1_mux), .D(mult1_un187_sum_1_CO3_1_RNO), .Y(
        mult1_un187_sum_1_CO3_0));
    SLE \buff_0[0]  (.D(\k[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_0_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_0[0]_net_1 ));
    CFG3 #( .INIT(8'h2E) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM[4]  (.A(
        \mult1_un159_sum_1_SUM[4] ), .B(
        \mult1_un159_sum_1_SUM_RNIM44K4[4] ), .C(
        \mult1_un159_sum_1_SUM[2] ), .Y(\mult1_un166_sum_1_SUM[4] ));
    CFG4 #( .INIT(16'h3A30) )  \i_lm_0[2]  (.A(\i_s[2] ), .B(N_144), 
        .C(\state[4]_net_1 ), .D(N_91), .Y(\i_lm[2] ));
    CFG2 #( .INIT(4'h9) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM_0[1]  (.A(
        \valu[5]_net_1 ), .B(\valu[6]_net_1 ), .Y(d_N_4_1));
    CFG4 #( .INIT(16'h3933) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_CO3_1_RNO  (.A(
        mult1_un180_sum_1_CO3_1), .B(\mult1_un180_sum_1_SUM_2[4] ), .C(
        mult1_un180_sum_1_CO3_a4), .D(mult1_un180_sum_1_CO3_0_0), .Y(
        mult1_un187_sum_1_CO3_1_RNO));
    CFG4 #( .INIT(16'h2AEA) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO_2  (.A(
        \mult1_un194_sum_1_SUM_1[4] ), .B(\mult1_un187_sum_1_SUM[1] ), 
        .C(\mult1_un187_sum_1_SUM[2] ), .D(d_N_2_0), .Y(d_N_11_mux));
    CFG2 #( .INIT(4'hD) )  \un1_angle[4]  (.A(\state[4]_net_1 ), .B(
        \k[5] ), .Y(\un1_angle[4]_net_1 ));
    CFG4 #( .INIT(16'hC0AF) )  \data_out_1_5_am[4]  (.A(\buff_5[5] ), 
        .B(\buff_4[5] ), .C(\i[2]_net_1 ), .D(
        \data_out_1_5_am_1_1[4]_net_1 ), .Y(\data_out_1_5_am[4]_net_1 )
        );
    CFG3 #( .INIT(8'hD8) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_CO2_1  (.A(
        un1_i1_mux), .B(\mult1_un180_sum_1_SUM[4] ), .C(
        \mult1_un180_sum_1_SUM[1] ), .Y(mult1_un187_sum_1_CO2));
    CFG4 #( .INIT(16'h24DB) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM[2]  (.A(
        \valu[10]_net_1 ), .B(\valu[11]_net_1 ), .C(
        \valu_RNI32OE1[13]_net_1 ), .D(\valu_RNILKIF_0[11]_net_1 ), .Y(
        \mult1_un159_sum_1_SUM[2] ));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM[4]  (.A(
        \valu_RNI32OE1[13]_net_1 ), .B(mult1_un159_sum_1_CO3), .C(
        \mult1_un159_sum_1_SUM_2_1[4] ), .Y(\mult1_un159_sum_1_SUM[4] )
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_23 (.A(VCC_net_1), .B(
        \i[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_22_net_1), .S(un1_i_cry_23_S_0), .Y(), .FCO(
        un1_i_cry_23_net_1));
    CFG4 #( .INIT(16'hAE2A) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO2_1  (.A(
        \mult1_un173_sum_1_SUM[1] ), .B(un1_i3_mux_0_0_i), .C(
        \valu[8]_net_1 ), .D(\valu[7]_net_1 ), .Y(
        mult1_un180_sum_1_CO2));
    SLE \data_out[1]  (.D(\data_out_1[1] ), .CLK(FCCC_0_GL0), .EN(
        data_out_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        time_sender_0_data_out_1));
    SLE \buff_0[2]  (.D(\k[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_0_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_0[2]_net_1 ));
    CFG4 #( .INIT(16'hFD10) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_CO3_1  (.A(
        \valu_RNI32OE1[13]_net_1 ), .B(un1_m5_i_0), .C(
        \valu_RNILKIF_0[11]_net_1 ), .D(\valu_RNICB5V[13]_net_1 ), .Y(
        mult1_un159_sum_1_CO3));
    SLE \buff_4[4]  (.D(\k[5] ), .CLK(FCCC_0_GL0), .EN(
        buff_4_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\buff_4[5] ));
    SLE \valu[7]  (.D(\un1_time1[7]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[7]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  buff_2_1_sqmuxa_1 (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(buff_2_1_sqmuxa_net_1), .D(\i[0]_net_1 ), .Y(
        buff_2_1_sqmuxa_1_net_1));
    CFG3 #( .INIT(8'h80) )  \state_ns_a2_0_a3[6]  (.A(
        \state_ns_i_0_a2_20[5]_net_1 ), .B(\state[2]_net_1 ), .C(
        \state_ns_i_0_a2_21[5]_net_1 ), .Y(\state_ns[6] ));
    SLE \buff_2[0]  (.D(\k[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_2_1_sqmuxa_1_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_2[0]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_bm[3]  (.A(\buff_2[3]_net_1 )
        , .B(\i[0]_net_1 ), .C(\buff_3[3]_net_1 ), .Y(
        \data_out_1_5_bm[3]_net_1 ));
    CFG4 #( .INIT(16'h5695) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_SUM[2]  (.A(
        \mult1_un173_sum_1_SUM[1] ), .B(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .C(\valu[8]_net_1 ), .D(
        \valu[7]_net_1 ), .Y(\mult1_un180_sum_1_SUM[2] ));
    SLE \buff_0[4]  (.D(\k[5] ), .CLK(FCCC_0_GL0), .EN(buff_0_1_sqmuxa)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\buff_0[5] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_21 (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_20_net_1), .S(un1_i_cry_21_S), .Y(), .FCO(
        un1_i_cry_21_net_1));
    CFG2 #( .INIT(4'h7) )  \state_ns_i_o2_0[1]  (.A(
        pulse_meash_0_new_ready), .B(\state[6]_net_1 ), .Y(N_91));
    SLE \valu[13]  (.D(\un1_time1[13]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[13]_net_1 ));
    CFG4 #( .INIT(16'hCEEE) )  \state_ns_i_0_a2_20_RNILRIH1[5]  (.A(
        \state[2]_net_1 ), .B(\un1_clk_inv_i_0_o3[0]_net_1 ), .C(
        \state_ns_i_0_a2_21[5]_net_1 ), .D(
        \state_ns_i_0_a2_20[5]_net_1 ), .Y(N_84_i_0));
    SLE \buff_5[1]  (.D(\k[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_5_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_5[1]_net_1 ));
    SLE \state[4]  (.D(\state[5]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\state[4]_net_1 ));
    CFG4 #( .INIT(16'hA2BA) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO2  (.A(
        \mult1_un208_sum_1_SUM[1] ), .B(
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] ), .C(\valu[2]_net_1 ), .D(
        \valu[3]_net_1 ), .Y(mult1_un215_sum_1_CO2));
    CFG4 #( .INIT(16'h2262) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM_RNITTTU_0[2]  (
        .A(\mult1_un166_sum_1_SUM[2] ), .B(mult1_un166_sum_1_CO3), .C(
        \valu[9]_net_1 ), .D(\valu[8]_net_1 ), .Y(un1_N_13_mux));
    CFG2 #( .INIT(4'hD) )  \state_ns_i_o2_0[3]  (.A(\state[3]_net_1 ), 
        .B(COREUART_0_TXRDY), .Y(N_90));
    CFG4 #( .INIT(16'h0020) )  buff_4_1_sqmuxa (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(buff_2_1_sqmuxa_net_1), .D(\i[0]_net_1 ), .Y(
        buff_4_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'h3237) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1  (.A(
        un1_m8_i_0), .B(d_i6_mux_1), .C(un1_N_7_0), .D(
        mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK), .Y(
        mult1_un201_sum_1_CO1));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[25]  (.A(\i_s[25]_net_1 ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[25] ));
    SLE \valu[3]  (.D(\un1_time1[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0_RNO_2  
        (.A(un1_i6_mux), .B(d_m12_0_a3_0), .Y(un1_N_10_mux));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM[1]  (.A(
        \valu[6]_net_1 ), .B(\mult1_un180_sum_1_SUM[4] ), .C(
        \valu[7]_net_1 ), .Y(\mult1_un187_sum_1_SUM[1] ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hAACF) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0  (.A(
        mult1_un201_sum_1_CO3_0_tz_s_0_RNO), .B(d_N_20), .C(d_N_19), 
        .D(un1_N_10_mux), .Y(mult1_un201_sum_1_CO3_0_tz_s_0));
    CFG2 #( .INIT(4'hB) )  \valu_RNILKIF[11]  (.A(\valu[12]_net_1 ), 
        .B(\valu[11]_net_1 ), .Y(un1_N_3_mux));
    SLE \buff_5[3]  (.D(\k[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_5_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_5[3]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  buff_3_1_sqmuxa (.A(\i[2]_net_1 ), .B(
        \i[1]_net_1 ), .C(buff_2_1_sqmuxa_net_1), .D(\i[0]_net_1 ), .Y(
        buff_3_1_sqmuxa_net_1));
    SLE \buff_0[1]  (.D(\k[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_0_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_0[1]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \un1_angle[1]  (.A(
        locator_control_0_angle1[1]), .B(\k[1]_net_1 ), .C(
        \state[4]_net_1 ), .Y(\un1_angle[1]_net_1 ));
    CFG4 #( .INIT(16'h05F3) )  \data_out_1_5_am_1_1[4]  (.A(
        \buff_1[5] ), .B(\buff_0[5] ), .C(\i[2]_net_1 ), .D(
        \i[0]_net_1 ), .Y(\data_out_1_5_am_1_1[4]_net_1 ));
    CFG3 #( .INIT(8'h2E) )  \un1_time1[9]  (.A(pulse_meash_0_tim[9]), 
        .B(\state[4]_net_1 ), .C(\mult1_un159_sum_1_SUM[4] ), .Y(
        \un1_time1[9]_net_1 ));
    SLE \i[23]  (.D(\i_lm[23] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[23]_net_1 ));
    CFG4 #( .INIT(16'hD44D) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_RNI6RET  (.A(
        \valu[2]_net_1 ), .B(\valu[1]_net_1 ), .C(
        mult1_un215_sum_1_CO3), .D(\mult1_un215_sum_1_SUM_0[4] ), .Y(
        mult1_un222_sum_1_CO1));
    CFG4 #( .INIT(16'hC3BE) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO3_2_0  (.A(
        \valu[7]_net_1 ), .B(\mult1_un166_sum_1_SUM[4] ), .C(
        \valu[9]_net_1 ), .D(\valu[8]_net_1 ), .Y(
        mult1_un180_sum_1_CO3_2_0));
    SLE \state[5]  (.D(N_85_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[5]_net_1 ));
    CFG4 #( .INIT(16'h5D75) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM_RNIM44K4[4]  (.A(
        un1_N_5_i_1), .B(\mult1_un159_sum_1_SUM[4] ), .C(
        \valu[10]_net_1 ), .D(\valu[9]_net_1 ), .Y(
        \mult1_un159_sum_1_SUM_RNIM44K4[4] ));
    SLE \buff_3[0]  (.D(\k[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_3_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_3[0]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  buff_0_1_sqmuxa_0_a2_0_a3 (.A(
        \i[0]_net_1 ), .B(\state[4]_net_1 ), .C(\i[1]_net_1 ), .D(
        \i[2]_net_1 ), .Y(buff_0_1_sqmuxa));
    ARI1 #( .INIT(20'h65500) )  \i_cry[23]  (.A(VCC_net_1), .B(
        \i[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[22]_net_1 ), .S(\i_s[23] ), .Y(), .FCO(
        \i_cry[23]_net_1 ));
    SLE \i[13]  (.D(\i_lm[13] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    CFG4 #( .INIT(16'hBEEB) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0_RNO_3  (.A(
        \valu[4]_net_1 ), .B(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), 
        .C(\mult1_un194_sum_1_SUM[1] ), .D(mult1_un201_sum_1_CO1), .Y(
        un1_N_8));
    CFG4 #( .INIT(16'hB000) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO_1  (.A(
        \valu[5]_net_1 ), .B(\valu[6]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[2] ), .D(\mult1_un187_sum_1_SUM[1] ), 
        .Y(un1_N_7_0));
    SLE \buff_1[1]  (.D(\un1_angle[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_2_i_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_1[1]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[15]  (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[14]_net_1 ), .S(\i_s[15] ), .Y(), .FCO(
        \i_cry[15]_net_1 ));
    CFG2 #( .INIT(4'h8) )  buff_2_1_sqmuxa (.A(\state[4]_net_1 ), .B(
        FCCC_0_LOCK), .Y(buff_2_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'hC693) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM_RNIQ5884[1]  (.A(
        \mult1_un166_sum_1_SUM[1] ), .B(un1_m8_1), .C(un1_N_13_mux), 
        .D(un1_i4_mux), .Y(\mult1_un166_sum_1_SUM_RNIQ5884[1] ));
    CFG2 #( .INIT(4'h7) )  \state_ns_i_o2[3]  (.A(un15_clklto2), .B(
        un15_clklto1), .Y(N_89));
    CFG3 #( .INIT(8'h28) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO_4  (.A(
        \valu[6]_net_1 ), .B(\mult1_un180_sum_1_SUM[4] ), .C(
        \valu[7]_net_1 ), .Y(d_N_12_0));
    CFG2 #( .INIT(4'h6) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM_RNIMGHHA[2]  (.A(
        un1_i2_mux), .B(un1_m6_1_0), .Y(
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_0_a2_16[5]  (.A(
        \i[15]_net_1 ), .B(\i[14]_net_1 ), .C(\i[11]_net_1 ), .D(
        \i[10]_net_1 ), .Y(\state_ns_i_0_a2_16[5]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  \i_8_iv_i_a2[2]  (.A(
        \state_ns_i_a2_17[3]_net_1 ), .B(\state_ns_i_a2_21[3]_net_1 ), 
        .C(un15_clklto2), .D(\state_ns_i_a2_16[3]_net_1 ), .Y(N_144));
    CFG3 #( .INIT(8'hF2) )  un1_rst_n_inv_2_i_0 (.A(FCCC_0_LOCK), .B(
        N_91), .C(N_104), .Y(un1_rst_n_inv_2_i_0_net_1));
    CFG4 #( .INIT(16'h1F10) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC3_0_RNO_0  (.A(
        d_N_10), .B(\mult1_un187_sum_1_SUM[1] ), .C(
        \mult1_un187_sum_1_SUM[4] ), .D(d_i5_mux), .Y(
        mult1_un201_sum_1_ANC3_0_RNO_0));
    SLE \k[4]  (.D(VCC_net_1), .CLK(FCCC_0_GL0), .EN(N_87_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\k[5] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[10]  (.A(\i_s[10] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[10] ));
    CFG4 #( .INIT(16'h9669) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO2_RNILDOT2  (.A(
        \mult1_un187_sum_1_SUM[2] ), .B(\mult1_un187_sum_1_SUM[4] ), 
        .C(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .D(
        mult1_un194_sum_1_CO2), .Y(\mult1_un201_sum_1_SUM_2[4] ));
    CFG3 #( .INIT(8'h57) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM_RNI6LH01[2]  (.A(
        \mult1_un187_sum_1_SUM[2] ), .B(d_m2_3_0), .C(
        \mult1_un187_sum_1_SUM[1] ), .Y(un1_m9_1));
    SLE \data_out[2]  (.D(\data_out_1[2] ), .CLK(FCCC_0_GL0), .EN(
        data_out_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        time_sender_0_data_out_2));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_s_1_323 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(un1_i_s_1_323_FCO));
    SLE \i[17]  (.D(\i_lm[17] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[17]_net_1 ));
    CFG4 #( .INIT(16'h1ED2) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42  
        (.A(un1_m9_1), .B(mult1_un187_sum_1_CO3_1_RNIDREF), .C(
        \mult1_un194_sum_1_SUM_1[4] ), .D(mult1_un194_sum_1_CO3_0_tz), 
        .Y(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42));
    CFG4 #( .INIT(16'h7340) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_ANC3_0_1  (.A(
        mult1_un194_sum_1_ANC3_0_1_1), .B(\mult1_un187_sum_1_SUM[4] ), 
        .C(\mult1_un187_sum_1_SUM[2] ), .D(mult1_un194_sum_1_CO3_0_tz), 
        .Y(mult1_un194_sum_1_ANC3_0_1));
    CFG4 #( .INIT(16'hECFE) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO2_0_tz  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .B(
        \mult1_un194_sum_1_SUM[1] ), .C(\valu[4]_net_1 ), .D(
        \valu[5]_net_1 ), .Y(mult1_un201_sum_1_CO2_0_tz));
    SLE \buff_5[0]  (.D(\k[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_5_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_5[0]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  wen_RNO_0 (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .C(\state[2]_net_1 ), .Y(N_445_i_0));
    CFG4 #( .INIT(16'hBA32) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO_0  (.A(
        \valu[5]_net_1 ), .B(\valu[4]_net_1 ), .C(d_N_11_mux), .D(
        d_N_13_mux), .Y(d_i6_mux_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_7 (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_6_net_1), .S(un1_i_cry_7_S_0), .Y(), .FCO(
        un1_i_cry_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_4 (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_3_net_1), .S(un1_i_cry_4_S_0), .Y(), .FCO(
        un1_i_cry_4_net_1));
    SLE \k[2]  (.D(\un24_k_v[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_87_i_0), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\k[2]_net_1 ));
    CFG3 #( .INIT(8'h42) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM_RNIEMCS[1]  (.A(
        \valu[9]_net_1 ), .B(\mult1_un159_sum_1_SUM[1] ), .C(
        \valu[10]_net_1 ), .Y(un1_m8_1_1));
    SLE \valu[9]  (.D(\un1_time1[9]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[9]_net_1 ));
    CFG4 #( .INIT(16'hC0AF) )  \data_out_1_5_am[3]  (.A(
        \buff_5[3]_net_1 ), .B(\buff_4[3]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\data_out_1_5_am_1_1[3]_net_1 ), .Y(
        \data_out_1_5_am[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \valu_RNIRVUG[5]  (.A(\valu[5]_net_1 ), .B(
        \valu[6]_net_1 ), .Y(d_m2_3_0));
    CFG4 #( .INIT(16'hFD40) )  
        \un1_k_if_generate_plus.mult1_un222_sum_1_CO3_1  (.A(
        \mult1_un215_sum_1_SUM[4] ), .B(mult1_un222_sum_1_CO1), .C(
        \mult1_un215_sum_1_SUM[1] ), .D(\mult1_un215_sum_1_SUM[2] ), 
        .Y(mult1_un222_sum_1_CO3));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_12[3]  (.A(
        un1_i_cry_3_S_0), .B(un1_i_cry_4_S_0), .C(un1_i_cry_5_S_0), .D(
        un1_i_cry_6_S_0), .Y(\state_ns_i_a2_12[3]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[17]  (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[16]_net_1 ), .S(\i_s[17] ), .Y(), .FCO(
        \i_cry[17]_net_1 ));
    CFG3 #( .INIT(8'h4C) )  \state_RNO[1]  (.A(
        \state_ns_i_0_a2_20[5]_net_1 ), .B(\state[2]_net_1 ), .C(
        \state_ns_i_0_a2_21[5]_net_1 ), .Y(N_84_tz_i));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[18]  (.A(\i_s[18] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[18] ));
    SLE \valu[4]  (.D(\un1_time1[4]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[4]_net_1 ));
    SLE \i[9]  (.D(\i_lm[9] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un208_sum_1_SUM[1]  (.A(
        \valu[4]_net_1 ), .B(\valu[3]_net_1 ), .C(
        mult1_un201_sum_1_CO3), .D(\mult1_un201_sum_1_SUM_2[4] ), .Y(
        \mult1_un208_sum_1_SUM[1] ));
    CFG4 #( .INIT(16'h4666) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO2_0_d_0_RNO  (.A(
        \valu[5]_net_1 ), .B(\valu[6]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[2] ), .D(\mult1_un187_sum_1_SUM[1] ), 
        .Y(un1_N_7_mux_0));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_8 (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_7_net_1), .S(un1_i_cry_8_S), .Y(), .FCO(
        un1_i_cry_8_net_1));
    SLE \valu[5]  (.D(\un1_time1[5]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[5]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_0_a2_12[5]  (.A(
        \i[23]_net_1 ), .B(\i[22]_net_1 ), .C(\i[20]_net_1 ), .D(
        \i[19]_net_1 ), .Y(\state_ns_i_0_a2_12[5]_net_1 ));
    CFG4 #( .INIT(16'h7800) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0_RNO_0  (.A(
        \mult1_un201_sum_1_SUM[2] ), .B(\mult1_un201_sum_1_SUM[4] ), 
        .C(un1_N_5_mux), .D(un1_m7_3_0), .Y(un1_i5_mux_0));
    CFG2 #( .INIT(4'hE) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_0  (.A(
        mult1_un201_sum_1_CO3_0_0_1), .B(mult1_un201_sum_1_CO3_0_d), 
        .Y(mult1_un201_sum_1_CO3));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_16[3]  (.A(
        un1_i_cry_18_S_0), .B(un1_i_cry_19_S_0), .C(un1_i_cry_20_S), 
        .D(un1_i_cry_21_S), .Y(\state_ns_i_a2_16[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \buff_2[2]  (.D(\k[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_2_1_sqmuxa_1_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_2[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM[1]  (.A(
        mult1_un194_sum_1_ANC3_0_1), .B(\mult1_un201_sum_1_SUM_1[1] ), 
        .Y(N_3560_i));
    CFG3 #( .INIT(8'h40) )  \i_8_iv_i_a3[1]  (.A(un15_clklto2), .B(
        \state_ns_i_a2[3]_net_1 ), .C(un15_clklto1), .Y(N_95));
    SLE \valu[0]  (.D(\un1_time1[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_12 (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_11_net_1), .S(un1_i_cry_12_S_0), .Y(), .FCO(
        un1_i_cry_12_net_1));
    CFG4 #( .INIT(16'h444B) )  \valu_RNI32OE1_0[13]  (.A(
        \valu_RNINMIF[13]_net_1 ), .B(un1_N_3_mux), .C(
        \valu[13]_net_1 ), .D(\valu[12]_net_1 ), .Y(
        \mult1_un159_sum_1_SUM_2_1[4] ));
    CFG4 #( .INIT(16'h0012) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC3_0_RNO  (.A(
        \valu[4]_net_1 ), .B(\valu[6]_net_1 ), .C(\valu[5]_net_1 ), .D(
        \mult1_un187_sum_1_SUM[1] ), .Y(un1_m4_1_1));
    CFG4 #( .INIT(16'h3CE1) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0_RNO_2  (.A(
        mult1_un201_sum_1_CO2_0_tz), .B(mult1_un201_sum_1_ANC2), .C(
        \valu[3]_net_1 ), .D(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), 
        .Y(un1_m7_i_0_1));
    CFG4 #( .INIT(16'h5A33) )  
        \un1_k_if_generate_plus.mult1_un208_sum_1_CO2_1  (.A(
        \mult1_un201_sum_1_SUM_2[4] ), .B(N_3560_i), .C(
        mult1_un201_sum_1_CO3), .D(un1_i3_mux_0), .Y(
        mult1_un208_sum_1_CO2));
    CFG4 #( .INIT(16'hFE01) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_c_RNI45FP3  (
        .A(mult1_un201_sum_1_CO3_0_c), .B(mult1_un201_sum_1_CO3_0_d), 
        .C(mult1_un201_sum_1_ANC3), .D(\mult1_un201_sum_1_SUM_2[4] ), 
        .Y(mult1_un201_sum_1_CO3_0_c_RNI45FP3));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM_0_RNIIHPG[4]  (
        .A(\mult1_un180_sum_1_SUM[2] ), .B(\mult1_un180_sum_1_SUM[4] ), 
        .C(mult1_un187_sum_1_CO2), .D(\mult1_un187_sum_1_SUM_0[4] ), 
        .Y(d_m1_2_0));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_15[3]  (.A(
        un1_i_cry_25_net_1), .B(un1_i_cry_15_S_0), .C(un1_i_cry_16_S_0)
        , .D(un1_i_cry_17_S), .Y(\state_ns_i_a2_15[3]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \un24_k_v_1[1]  (.A(\valu[2]_net_1 ), 
        .B(\valu[1]_net_1 ), .C(mult1_un215_sum_1_CO3), .D(
        \mult1_un215_sum_1_SUM_0[4] ), .Y(\un24_k_v_1[1]_net_1 ));
    CFG4 #( .INIT(16'h7080) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0_RNO_0  
        (.A(\mult1_un187_sum_1_SUM[2] ), .B(\mult1_un187_sum_1_SUM[4] )
        , .C(d_m12_0_a3_0), .D(\mult1_un194_sum_1_SUM_1[4] ), .Y(
        d_N_20));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_ns[1]  (.A(
        \data_out_1_5_am[1]_net_1 ), .B(\i[1]_net_1 ), .C(
        \data_out_1_5_bm[1]_net_1 ), .Y(\data_out_1[1] ));
    CFG4 #( .INIT(16'h572A) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC3_0_RNO_1  (.A(
        \valu[6]_net_1 ), .B(\valu[4]_net_1 ), .C(
        \mult1_un194_sum_1_SUM_1[4] ), .D(\valu[5]_net_1 ), .Y(d_N_10));
    CFG4 #( .INIT(16'hD2B4) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM_0_0[3]  (.A(
        \valu[3]_net_1 ), .B(\valu[4]_net_1 ), .C(N_3560_i), .D(
        \mult1_un201_sum_1_SUM[4] ), .Y(\mult1_un215_sum_1_SUM_0[3] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_5 (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_4_net_1), .S(un1_i_cry_5_S_0), .Y(), .FCO(
        un1_i_cry_5_net_1));
    CFG4 #( .INIT(16'h05F3) )  \data_out_1_5_am_1_1[0]  (.A(
        \buff_1[0]_net_1 ), .B(\buff_0[0]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\i[0]_net_1 ), .Y(\data_out_1_5_am_1_1[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_10 (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_9_net_1), .S(un1_i_cry_10_S_0), .Y(), .FCO(
        un1_i_cry_10_net_1));
    CFG4 #( .INIT(16'h99BD) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM_RNISQFG7[2]  (.A(
        \mult1_un201_sum_1_SUM[2] ), .B(
        mult1_un201_sum_1_CO3_0_c_RNI45FP3), .C(N_3560_i), .D(
        un1_i3_mux_0), .Y(un1_i2_mux));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un222_sum_1_SUM_0[4]  (.A(
        mult1_un215_sum_1_CO2), .B(\mult1_un215_sum_1_SUM[4] ), .C(
        \mult1_un215_sum_1_SUM_1[3] ), .Y(\mult1_un222_sum_1_SUM_0[4] )
        );
    CFG3 #( .INIT(8'hF8) )  \un1_clk_inv_i_0_o3[0]  (.A(
        \state[6]_net_1 ), .B(pulse_meash_0_new_ready), .C(
        \state[4]_net_1 ), .Y(\un1_clk_inv_i_0_o3[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  wen_RNIIK85 (.A(LED_3_c), .Y(LED_3_c_i_0));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_SUM[1]  (.A(
        \valu[8]_net_1 ), .B(\valu[7]_net_1 ), .C(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .Y(
        \mult1_un180_sum_1_SUM[1] ));
    CFG4 #( .INIT(16'h4DD4) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO1  (.A(
        \valu[3]_net_1 ), .B(\valu[2]_net_1 ), .C(un1_i2_mux), .D(
        un1_m6_1_0), .Y(mult1_un215_sum_1_CO1));
    CFG3 #( .INIT(8'h2E) )  \un1_time1[10]  (.A(pulse_meash_0_tim[10]), 
        .B(\state[4]_net_1 ), .C(\valu_RNI32OE1[13]_net_1 ), .Y(
        \un1_time1[10]_net_1 ));
    CFG4 #( .INIT(16'hFE88) )  
        \un1_k_if_generate_plus.mult1_un173_sum_1_CO2  (.A(
        mult1_un173_sum_1_CO1_0), .B(\mult1_un166_sum_1_SUM[4] ), .C(
        \valu[8]_net_1 ), .D(\mult1_un166_sum_1_SUM[1] ), .Y(
        mult1_un173_sum_1_CO2));
    CFG2 #( .INIT(4'h8) )  \state_RNO[2]  (.A(\state[3]_net_1 ), .B(
        COREUART_0_TXRDY), .Y(N_431_i_0));
    ARI1 #( .INIT(20'h45500) )  \i_s[25]  (.A(VCC_net_1), .B(
        \i[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[24]_net_1 ), .S(\i_s[25]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_6 (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_5_net_1), .S(un1_i_cry_6_S_0), .Y(), .FCO(
        un1_i_cry_6_net_1));
    ARI1 #( .INIT(20'h65500) )  \i_cry[11]  (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[10]_net_1 ), .S(\i_s[11] ), .Y(), .FCO(
        \i_cry[11]_net_1 ));
    SLE \buff_4[2]  (.D(\k[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_4_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_4[2]_net_1 ));
    CFG4 #( .INIT(16'hEEAE) )  
        \un1_k_if_generate_plus.mult1_un173_sum_1_SUM_RNIQIB05[2]  (.A(
        \mult1_un173_sum_1_SUM[2] ), .B(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .C(\valu[8]_net_1 ), .D(
        \valu[7]_net_1 ), .Y(mult1_un180_sum_1_CO3_1));
    CFG2 #( .INIT(4'h1) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO3_a4  (.A(
        \mult1_un173_sum_1_SUM[1] ), .B(\mult1_un173_sum_1_SUM[2] ), 
        .Y(mult1_un180_sum_1_CO3_a4));
    SLE \i[25]  (.D(\i_lm[25] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[25]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_1 (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_s_1_323_FCO), .S(un15_clklto1), .Y(), .FCO(
        un1_i_cry_1_net_1));
    SLE \k[3]  (.D(\SUM[3] ), .CLK(FCCC_0_GL0), .EN(N_87_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\k[3]_net_1 ));
    SLE \k[0]  (.D(\valu[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(N_87_i_0), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\k[0]_net_1 ));
    SLE \buff_3[3]  (.D(\k[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_3_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_3[3]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[24]  (.A(VCC_net_1), .B(
        \i[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[23]_net_1 ), .S(\i_s[24] ), .Y(), .FCO(
        \i_cry[24]_net_1 ));
    CFG4 #( .INIT(16'h2409) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0_RNO  (.A(
        \valu[3]_net_1 ), .B(\valu[4]_net_1 ), .C(N_3560_i), .D(
        \mult1_un201_sum_1_SUM[4] ), .Y(mult1_un215_sum_1_CO3_0_RNO));
    CFG2 #( .INIT(4'hE) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO3_2  (.A(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .B(
        mult1_un180_sum_1_CO3_2_0), .Y(mult1_un180_sum_1_CO3_0_0));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[19]  (.A(\i_s[19] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[19] ));
    SLE \i[15]  (.D(\i_lm[15] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[15]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[3]  (.A(\i_s[3] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[3] ));
    CFG4 #( .INIT(16'h1E5A) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM[4]  (.A(
        mult1_un187_sum_1_CO3_0), .B(\mult1_un180_sum_1_SUM[2] ), .C(
        \mult1_un187_sum_1_SUM_0[4] ), .D(mult1_un187_sum_1_CO2), .Y(
        \mult1_un187_sum_1_SUM[4] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[16]  (.A(\i_s[16] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[16] ));
    SLE wen (.D(N_139_i_0), .CLK(FCCC_0_GL0), .EN(N_445_i_0), .ALn(
        FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(LED_3_c));
    CFG4 #( .INIT(16'h05F3) )  \data_out_1_5_am_1_1[2]  (.A(
        \buff_1[2]_net_1 ), .B(\buff_0[2]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\i[0]_net_1 ), .Y(\data_out_1_5_am_1_1[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[20]  (.A(\i_s[20] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[20] ));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un1_sum_1.SUM_1[3]  (.A(
        \mult1_un215_sum_1_SUM_0[4] ), .B(\mult1_un215_sum_1_SUM[1] ), 
        .C(mult1_un222_sum_1_CO1), .D(mult1_un215_sum_1_CO3), .Y(
        \SUM_1[3] ));
    CFG2 #( .INIT(4'hE) )  wen_RNO (.A(\state[1]_net_1 ), .B(
        \state[0]_net_1 ), .Y(N_139_i_0));
    CFG2 #( .INIT(4'h6) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO2_1_RNO_0  (.A(
        un1_m8_1), .B(\valu[7]_net_1 ), .Y(un1_m2_5_0));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un1_sum_1.SUM[3]  (.A(\SUM_1[3] )
        , .B(mult1_un222_sum_1_CO3), .C(CO2), .D(
        \mult1_un222_sum_1_SUM_0[4] ), .Y(\SUM[3] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7] ), .Y(), .FCO(\i_cry[7]_net_1 ));
    CFG2 #( .INIT(4'h9) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0_RNO_3  (.A(
        \mult1_un194_sum_1_SUM[2] ), .B(\valu[3]_net_1 ), .Y(
        mult1_un215_sum_1_CO3_0_RNO_3));
    CFG4 #( .INIT(16'hB888) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO2_0_d_0_RNO_0  (.A(
        d_N_11_mux_0), .B(\mult1_un187_sum_1_SUM[4] ), .C(d_m2_3_0), 
        .D(\mult1_un194_sum_1_SUM_1[4] ), .Y(
        mult1_un201_sum_1_CO2_0_d_0_RNO_0));
    SLE \i[22]  (.D(\i_lm[22] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[22]_net_1 ));
    CFG4 #( .INIT(16'hC99C) )  \un24_k_v[1]  (.A(\valu[1]_net_1 ), .B(
        \un24_k_v_1[1]_net_1 ), .C(\mult1_un222_sum_1_SUM_0[4] ), .D(
        mult1_un222_sum_1_CO3), .Y(\un24_k_v[1]_net_1 ));
    CFG3 #( .INIT(8'h18) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_CO3_1_RNO  (.A(
        \valu[10]_net_1 ), .B(\valu_RNICB5V[13]_net_1 ), .C(
        \valu[11]_net_1 ), .Y(un1_m5_i_0));
    ARI1 #( .INIT(20'h65500) )  \i_cry[12]  (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[11]_net_1 ), .S(\i_s[12] ), .Y(), .FCO(
        \i_cry[12]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \un1_time1[4]  (.A(pulse_meash_0_tim[4]), 
        .B(\state[4]_net_1 ), .C(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42)
        , .Y(\un1_time1[4]_net_1 ));
    CFG4 #( .INIT(16'h1E4B) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM_1[4]  (.A(
        un1_i1_mux), .B(\mult1_un180_sum_1_SUM[4] ), .C(
        \mult1_un180_sum_1_SUM[2] ), .D(\mult1_un180_sum_1_SUM[1] ), 
        .Y(\mult1_un194_sum_1_SUM_1[4] ));
    CFG4 #( .INIT(16'h24DB) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM[2]  (.A(
        \valu[5]_net_1 ), .B(\valu[6]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[4] ), .D(\mult1_un187_sum_1_SUM[1] ), 
        .Y(\mult1_un194_sum_1_SUM[2] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[6]  (.A(\i_s[6] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[6] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[18]  (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[17]_net_1 ), .S(\i_s[18] ), .Y(), .FCO(
        \i_cry[18]_net_1 ));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM_1[3]  (.A(
        \mult1_un215_sum_1_SUM_0[3] ), .B(un1_m6_1_0), .C(un1_i2_mux), 
        .Y(\mult1_un215_sum_1_SUM_1[3] ));
    CFG4 #( .INIT(16'h66C9) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0_RNO_1  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .B(
        mult1_un215_sum_1_CO3_0_RNO_3), .C(mult1_un201_sum_1_CO2_0_tz), 
        .D(mult1_un201_sum_1_ANC2), .Y(un1_N_5_mux));
    SLE \i[2]  (.D(\i_lm[2] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \valu_RNINMIF[13]  (.A(\valu[12]_net_1 ), 
        .B(\valu[13]_net_1 ), .Y(\valu_RNINMIF[13]_net_1 ));
    CFG3 #( .INIT(8'h56) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM[4]  (.A(
        \mult1_un201_sum_1_SUM_2[4] ), .B(mult1_un201_sum_1_CO3_0_d), 
        .C(mult1_un201_sum_1_CO3_0_0_1), .Y(\mult1_un201_sum_1_SUM[4] )
        );
    CFG4 #( .INIT(16'h9669) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_SUM_2[4]  (.A(
        \mult1_un166_sum_1_SUM[4] ), .B(\mult1_un166_sum_1_SUM[2] ), 
        .C(\mult1_un166_sum_1_SUM_RNIQ5884[1] ), .D(
        mult1_un173_sum_1_CO2), .Y(\mult1_un180_sum_1_SUM_2[4] ));
    SLE \i[12]  (.D(\i_lm[12] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_15 (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_14_net_1), .S(un1_i_cry_15_S_0), .Y(), .FCO(
        un1_i_cry_15_net_1));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_ns[3]  (.A(
        \data_out_1_5_am[3]_net_1 ), .B(\i[1]_net_1 ), .C(
        \data_out_1_5_bm[3]_net_1 ), .Y(\data_out_1[3] ));
    SLE \valu[8]  (.D(\un1_time1[8]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[8]_net_1 ));
    CFG4 #( .INIT(16'hC963) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_CO2_1_RNO  (.A(
        \mult1_un166_sum_1_SUM[1] ), .B(un1_m2_5_0), .C(un1_i4_mux), 
        .D(un1_N_13_mux), .Y(un1_i3_mux_0_0_i));
    CFG3 #( .INIT(8'h80) )  \state_ns_i_a2[3]  (.A(
        \state_ns_i_a2_16[3]_net_1 ), .B(\state_ns_i_a2_17[3]_net_1 ), 
        .C(\state_ns_i_a2_21[3]_net_1 ), .Y(\state_ns_i_a2[3]_net_1 ));
    CFG4 #( .INIT(16'hE1A5) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_CO3_1_RNIDREF  (.A(
        mult1_un187_sum_1_CO3_0), .B(\mult1_un180_sum_1_SUM[2] ), .C(
        \mult1_un187_sum_1_SUM_0[4] ), .D(mult1_un187_sum_1_CO2), .Y(
        mult1_un187_sum_1_CO3_1_RNIDREF));
    CFG4 #( .INIT(16'hFB20) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO2  (.A(
        \valu[5]_net_1 ), .B(\valu[6]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[4] ), .D(\mult1_un187_sum_1_SUM[1] ), 
        .Y(mult1_un194_sum_1_CO2));
    CFG4 #( .INIT(16'hCACF) )  \i_lm_0[1]  (.A(\i_s[1] ), .B(N_95), .C(
        \state[4]_net_1 ), .D(N_91), .Y(\i_lm[1] ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_bm[1]  (.A(\buff_2[1]_net_1 )
        , .B(\i[0]_net_1 ), .C(\buff_3[1]_net_1 ), .Y(
        \data_out_1_5_bm[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \un1_time1[13]  (.A(\state[4]_net_1 ), .B(
        pulse_meash_0_tim[13]), .Y(\un1_time1[13]_net_1 ));
    SLE \buff_4[0]  (.D(\k[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_4_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_4[0]_net_1 ));
    CFG4 #( .INIT(16'hE44E) )  \un1_time1[0]  (.A(\state[4]_net_1 ), 
        .B(pulse_meash_0_tim[0]), .C(mult1_un222_sum_1_CO3), .D(
        \mult1_un222_sum_1_SUM_0[4] ), .Y(\un1_time1[0]_net_1 ));
    CFG4 #( .INIT(16'h9996) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0_RNO  (.A(
        \valu[4]_net_1 ), .B(\mult1_un201_sum_1_SUM_2[4] ), .C(
        mult1_un201_sum_1_CO3_0_d), .D(mult1_un201_sum_1_CO3_0_0_1), 
        .Y(un1_N_7_i));
    CFG4 #( .INIT(16'h8976) )  
        \un1_k_if_generate_plus.mult1_un173_sum_1_SUM[2]  (.A(
        mult1_un173_sum_1_CO1_0), .B(\mult1_un166_sum_1_SUM[4] ), .C(
        \valu[8]_net_1 ), .D(\mult1_un166_sum_1_SUM[1] ), .Y(
        \mult1_un173_sum_1_SUM[2] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[12]  (.A(\i_s[12] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[12] ));
    SLE \buff_1[4]  (.D(\un1_angle[4]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_2_i_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_1[5] ));
    CFG4 #( .INIT(16'h5177) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM_RNI3FKB4[2]  (.A(
        \mult1_un159_sum_1_SUM[2] ), .B(
        mult1_un159_sum_1_CO3_1_RNI1HJB3), .C(\valu[10]_net_1 ), .D(
        \mult1_un159_sum_1_SUM[1] ), .Y(un1_N_5_1));
    SLE \i[20]  (.D(\i_lm[20] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[20]_net_1 ));
    SLE \data_out[3]  (.D(\data_out_1[3] ), .CLK(FCCC_0_GL0), .EN(
        data_out_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        time_sender_0_data_out_3));
    CFG4 #( .INIT(16'h0C20) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC3_0_RNO_2  (.A(
        \valu[4]_net_1 ), .B(\valu[6]_net_1 ), .C(\valu[5]_net_1 ), .D(
        \mult1_un187_sum_1_SUM[1] ), .Y(d_i5_mux));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_9 (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_8_net_1), .S(un1_i_cry_9_S_0), .Y(), .FCO(
        un1_i_cry_9_net_1));
    CFG4 #( .INIT(16'h05F3) )  \data_out_1_5_am_1_1[3]  (.A(
        \buff_1[3]_net_1 ), .B(\buff_0[3]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\i[0]_net_1 ), .Y(\data_out_1_5_am_1_1[3]_net_1 ));
    CFG4 #( .INIT(16'hC13E) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_SUM_RNIQL113[2]  (.A(
        mult1_un201_sum_1_CO2_0_tz), .B(mult1_un201_sum_1_ANC2), .C(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .D(
        \mult1_un194_sum_1_SUM[2] ), .Y(un1_m6_1_0));
    SLE \state[3]  (.D(N_10_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[11]  (.A(\i_s[11] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[11] ));
    CFG4 #( .INIT(16'h781E) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM[3]  (.A(
        mult1_un215_sum_1_CO1), .B(\mult1_un208_sum_1_SUM[1] ), .C(
        \mult1_un215_sum_1_SUM_1[3] ), .D(
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] ), .Y(
        \mult1_un215_sum_1_SUM[3] ));
    CFG3 #( .INIT(8'h80) )  data_out_0_sqmuxa_0_a3 (.A(FCCC_0_LOCK), 
        .B(COREUART_0_TXRDY), .C(\state[3]_net_1 ), .Y(
        data_out_0_sqmuxa));
    CFG2 #( .INIT(4'h4) )  \valu_RNO[11]  (.A(\state[4]_net_1 ), .B(
        pulse_meash_0_tim[11]), .Y(\valu_RNO[11]_net_1 ));
    SLE \valu[11]  (.D(\valu_RNO[11]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[11]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_18 (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_17_net_1), .S(un1_i_cry_18_S_0), .Y(), .FCO(
        un1_i_cry_18_net_1));
    SLE \i[10]  (.D(\i_lm[10] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    CFG2 #( .INIT(4'h6) )  
        \un1_k_if_generate_plus.mult1_un180_sum_1_SUM_0[3]  (.A(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .B(
        \mult1_un173_sum_1_SUM[2] ), .Y(\mult1_un180_sum_1_SUM_0[3] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_14 (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_13_net_1), .S(un1_i_cry_14_S_0), .Y(), .FCO(
        un1_i_cry_14_net_1));
    CFG4 #( .INIT(16'h0208) )  
        \un1_k_if_generate_plus.mult1_un1_sum_1.ANC2_0  (.A(ANC2_m3), 
        .B(\mult1_un215_sum_1_SUM[4] ), .C(\valu[1]_net_1 ), .D(
        \valu[2]_net_1 ), .Y(CO2));
    SLE \i[6]  (.D(\i_lm[6] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_bm[2]  (.A(\buff_2[2]_net_1 )
        , .B(\i[0]_net_1 ), .C(\buff_3[2]_net_1 ), .Y(
        \data_out_1_5_bm[2]_net_1 ));
    CFG4 #( .INIT(16'h7080) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO2_0_d_0_RNO_1  (.A(
        \mult1_un187_sum_1_SUM[1] ), .B(\mult1_un187_sum_1_SUM[2] ), 
        .C(d_N_4_1), .D(\mult1_un194_sum_1_SUM_1[4] ), .Y(d_N_11_mux_0)
        );
    ARI1 #( .INIT(20'h65500) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[0]_net_1 ), .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \un1_angle[0]  (.A(
        locator_control_0_angle1[0]), .B(\k[0]_net_1 ), .C(
        \state[4]_net_1 ), .Y(\un1_angle[0]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_lm[4] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[10]  (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[9]_net_1 ), .S(\i_s[10] ), .Y(), .FCO(\i_cry[10]_net_1 )
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_17 (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_16_net_1), .S(un1_i_cry_17_S), .Y(), .FCO(
        un1_i_cry_17_net_1));
    ARI1 #( .INIT(20'h65500) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    SLE \buff_3[4]  (.D(\k[5] ), .CLK(FCCC_0_GL0), .EN(
        buff_3_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\buff_3[5] ));
    CFG3 #( .INIT(8'hE2) )  \un1_time1[8]  (.A(pulse_meash_0_tim[8]), 
        .B(\state[4]_net_1 ), .C(mult1_un166_sum_1_CO3), .Y(
        \un1_time1[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_16 (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_15_net_1), .S(un1_i_cry_16_S_0), .Y(), .FCO(
        un1_i_cry_16_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_22 (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_21_net_1), .S(un1_i_cry_22_S_0), .Y(), .FCO(
        un1_i_cry_22_net_1));
    CFG4 #( .INIT(16'hF0F4) )  \state_ns_0[0]  (.A(
        pulse_meash_0_new_ready), .B(\state_ns_0_a3_3[0]_net_1 ), .C(
        \state[0]_net_1 ), .D(\state[4]_net_1 ), .Y(\state_ns[0] ));
    CFG4 #( .INIT(16'h7233) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_1), .B(
        mult1_un194_sum_1_CO3_0_tz_0_RNO), .C(\valu[5]_net_1 ), .D(
        \mult1_un180_sum_1_SUM[1] ), .Y(mult1_un194_sum_1_CO3_0_tz));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[8]  (.A(\i_s[8] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[8] ));
    SLE \i[19]  (.D(\i_lm[19] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[19]_net_1 ));
    CFG4 #( .INIT(16'h24DB) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM[2]  (.A(
        \valu[6]_net_1 ), .B(\valu[7]_net_1 ), .C(
        \mult1_un180_sum_1_SUM[4] ), .D(\mult1_un180_sum_1_SUM[1] ), 
        .Y(\mult1_un187_sum_1_SUM[2] ));
    CFG4 #( .INIT(16'h336C) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_CO3_1_RNI8N0S  (.A(
        mult1_un187_sum_1_CO2), .B(d_m1_2_0), .C(
        \mult1_un180_sum_1_SUM[2] ), .D(mult1_un187_sum_1_CO3_0), .Y(
        d_N_2_0));
    SLE \data_out[4]  (.D(\data_out_1[5] ), .CLK(FCCC_0_GL0), .EN(
        data_out_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        time_sender_0_data_out_5));
    SLE \buff_1[3]  (.D(\un1_angle[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_2_i_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_1[3]_net_1 ));
    CFG4 #( .INIT(16'h4EE4) )  \un1_time1[2]  (.A(\state[4]_net_1 ), 
        .B(pulse_meash_0_tim[2]), .C(un1_i2_mux), .D(un1_m6_1_0), .Y(
        \un1_time1[2]_net_1 ));
    CFG3 #( .INIT(8'h2E) )  \un1_time1[6]  (.A(pulse_meash_0_tim[6]), 
        .B(\state[4]_net_1 ), .C(\mult1_un180_sum_1_SUM[4] ), .Y(
        \un1_time1[6]_net_1 ));
    SLE \buff_2[1]  (.D(\k[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_2_1_sqmuxa_1_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_2[1]_net_1 ));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM[1]  (.A(
        \valu[9]_net_1 ), .B(\mult1_un159_sum_1_SUM[4] ), .C(
        \valu[10]_net_1 ), .Y(\mult1_un166_sum_1_SUM[1] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_20 (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_19_net_1), .S(un1_i_cry_20_S), .Y(), .FCO(
        un1_i_cry_20_net_1));
    CFG4 #( .INIT(16'h5965) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM[2]  (.A(
        \mult1_un208_sum_1_SUM[1] ), .B(
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] ), .C(\valu[2]_net_1 ), .D(
        \valu[3]_net_1 ), .Y(\mult1_un215_sum_1_SUM[2] ));
    CFG4 #( .INIT(16'h6669) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM_0_0[4]  (.A(
        \mult1_un201_sum_1_SUM[2] ), .B(\mult1_un201_sum_1_SUM_2[4] ), 
        .C(mult1_un201_sum_1_CO3_0_0_1), .D(mult1_un201_sum_1_CO3_0_d), 
        .Y(\mult1_un215_sum_1_SUM_0_0[4] ));
    SLE \buff_2[3]  (.D(\k[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_2_1_sqmuxa_1_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_2[3]_net_1 ));
    CFG4 #( .INIT(16'h1441) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0_RNO_2  (.A(
        N_3560_i), .B(\valu[4]_net_1 ), .C(mult1_un201_sum_1_CO3), .D(
        \mult1_un201_sum_1_SUM_2[4] ), .Y(un1_m7_3_0));
    CFG4 #( .INIT(16'hF4B0) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC3_0  (.A(
        \mult1_un187_sum_1_SUM[4] ), .B(un1_m4_1_1), .C(
        mult1_un201_sum_1_ANC3_0_RNO_0), .D(
        mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK), .Y(
        mult1_un201_sum_1_ANC3));
    CFG4 #( .INIT(16'hB54A) )  
        \un1_k_if_generate_plus.mult1_un1_sum_1.ANC2_m3  (.A(
        \valu[2]_net_1 ), .B(\mult1_un215_sum_1_SUM[1] ), .C(
        \mult1_un215_sum_1_SUM[2] ), .D(\mult1_un215_sum_1_SUM[3] ), 
        .Y(ANC2_m3));
    CFG4 #( .INIT(16'hD555) )  \state_RNO[5]  (.A(N_91), .B(
        \state[4]_net_1 ), .C(\state_ns_i_a2[3]_net_1 ), .D(N_89), .Y(
        N_85_i_0));
    SLE \buff_3[2]  (.D(\k[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_3_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_3[2]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \valu_RNILKIF_0[11]  (.A(\valu[12]_net_1 ), 
        .B(\valu[11]_net_1 ), .Y(\valu_RNILKIF_0[11]_net_1 ));
    CFG4 #( .INIT(16'h4920) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0_RNO  (.A(
        \valu[6]_net_1 ), .B(\valu[7]_net_1 ), .C(
        \mult1_un180_sum_1_SUM[4] ), .D(\mult1_un180_sum_1_SUM[1] ), 
        .Y(mult1_un194_sum_1_CO3_0_tz_0_RNO));
    SLE \i[24]  (.D(\i_lm[24] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[24]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_2 (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_1_net_1), .S(un15_clklto2), .Y(), .FCO(
        un1_i_cry_2_net_1));
    CFG4 #( .INIT(16'hC0AF) )  \data_out_1_5_am[1]  (.A(
        \buff_5[1]_net_1 ), .B(\buff_4[1]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\data_out_1_5_am_1_1[1]_net_1 ), .Y(
        \data_out_1_5_am[1]_net_1 ));
    CFG4 #( .INIT(16'hE44E) )  \un1_time1[1]  (.A(\state[4]_net_1 ), 
        .B(pulse_meash_0_tim[1]), .C(mult1_un215_sum_1_CO3), .D(
        \mult1_un215_sum_1_SUM_0[4] ), .Y(\un1_time1[1]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[7]  (.A(\i_s[7] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[7] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[13]  (.A(\i_s[13] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[13] ));
    CFG3 #( .INIT(8'hD1) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_CO3_1  (.A(
        \mult1_un159_sum_1_SUM[4] ), .B(
        \mult1_un159_sum_1_SUM_RNIM44K4[4] ), .C(
        \mult1_un159_sum_1_SUM[2] ), .Y(mult1_un166_sum_1_CO3));
    CFG4 #( .INIT(16'h40C0) )  \i_8_iv_i_a3[0]  (.A(un15_clklto2), .B(
        \state_ns_i_a2[3]_net_1 ), .C(\i[0]_net_1 ), .D(un15_clklto1), 
        .Y(N_96));
    CFG4 #( .INIT(16'h9669) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_CO3_1_RNI5BNN3  (.A(
        \valu_RNI32OE1[13]_net_1 ), .B(\mult1_un159_sum_1_SUM_2_1[4] ), 
        .C(mult1_un159_sum_1_CO3), .D(\mult1_un159_sum_1_SUM[1] ), .Y(
        un1_N_5_i_1));
    SLE \i[14]  (.D(\i_lm[14] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    SLE \state[2]  (.D(N_431_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  un1_rst_n_inv_i_a3 (.A(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .B(FCCC_0_LOCK), .Y(
        un1_rst_n_inv_i_a3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_3 (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_2_net_1), .S(un1_i_cry_3_S_0), .Y(), .FCO(
        un1_i_cry_3_net_1));
    CFG4 #( .INIT(16'h444F) )  \valu_RNI32OE1[13]  (.A(
        \valu_RNINMIF[13]_net_1 ), .B(un1_N_3_mux), .C(
        \valu[13]_net_1 ), .D(\valu[12]_net_1 ), .Y(
        \valu_RNI32OE1[13]_net_1 ));
    CFG4 #( .INIT(16'hF4B0) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO2_0_d_0  (.A(
        \mult1_un187_sum_1_SUM[4] ), .B(un1_N_7_mux_0), .C(
        mult1_un201_sum_1_CO2_0_d_0_RNO_0), .D(
        mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK), .Y(
        mult1_un201_sum_1_CO2_0_d));
    CFG4 #( .INIT(16'h8000) )  \state_ns_i_a2_21[3]  (.A(
        \state_ns_i_a2_12[3]_net_1 ), .B(\state_ns_i_a2_13[3]_net_1 ), 
        .C(\state_ns_i_a2_14[3]_net_1 ), .D(
        \state_ns_i_a2_15[3]_net_1 ), .Y(\state_ns_i_a2_21[3]_net_1 ));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0_1_RNO  (
        .A(\mult1_un180_sum_1_SUM_0[3] ), .B(\valu[6]_net_1 ), .C(
        mult1_un180_sum_1_CO2), .Y(mult1_un194_sum_1_CO3_0_tz_0_1_RNO));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_CO3_1_RNI1HJB3  (.A(
        \valu_RNI32OE1[13]_net_1 ), .B(mult1_un159_sum_1_CO3), .C(
        \mult1_un159_sum_1_SUM_2_1[4] ), .Y(
        mult1_un159_sum_1_CO3_1_RNI1HJB3));
    SLE \state[1]  (.D(N_84_tz_i), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    CFG4 #( .INIT(16'hC0AF) )  \data_out_1_5_am[2]  (.A(
        \buff_5[2]_net_1 ), .B(\buff_4[2]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\data_out_1_5_am_1_1[2]_net_1 ), .Y(
        \data_out_1_5_am[2]_net_1 ));
    CFG2 #( .INIT(4'h9) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK  
        (.A(mult1_un194_sum_1_CO3_0_tz), .B(
        \mult1_un194_sum_1_SUM_1[4] ), .Y(
        mult1_un194_sum_1_CO3_0_tz_0_RNIBNRK));
    ARI1 #( .INIT(20'h65500) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[22]  (.A(\i_s[22] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[22] ));
    SLE \i[5]  (.D(\i_lm[5] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    CFG3 #( .INIT(8'hA8) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_c  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .B(
        mult1_un201_sum_1_CO2_0_d), .C(mult1_un201_sum_1_CO3_0_tz_s_0), 
        .Y(mult1_un201_sum_1_CO3_0_c));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[9]  (.A(\i_s[9] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[9] ));
    SLE \i[8]  (.D(\i_lm[8] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    SLE \buff_1[2]  (.D(\un1_angle[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_2_i_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_1[2]_net_1 ));
    SLE \buff_4[3]  (.D(\k[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_4_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_4[3]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \un1_angle[3]  (.A(
        locator_control_0_angle1[3]), .B(\k[3]_net_1 ), .C(
        \state[4]_net_1 ), .Y(\un1_angle[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[21]  (.A(\i_s[21] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[21] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[13]  (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[12]_net_1 ), .S(\i_s[13] ), .Y(), .FCO(
        \i_cry[13]_net_1 ));
    SLE \valu[6]  (.D(\un1_time1[6]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[6]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[5]  (.A(\i_s[5] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[5] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_25 (.A(VCC_net_1), .B(
        \i[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_24_net_1), .S(un1_i_cry_25_S_0), .Y(), .FCO(
        un1_i_cry_25_net_1));
    CFG4 #( .INIT(16'h00EF) )  \state_RNO[3]  (.A(\state[1]_net_1 ), 
        .B(\state[4]_net_1 ), .C(N_90), .D(N_93), .Y(N_10_i_0));
    CFG2 #( .INIT(4'h8) )  \state_RNI45AA[5]  (.A(FCCC_0_LOCK), .B(
        \state[5]_net_1 ), .Y(N_87_i_0));
    CFG4 #( .INIT(16'h14EB) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM_RNIU8O02[2]  (.A(
        un1_m8_1_1), .B(\mult1_un159_sum_1_SUM[4] ), .C(
        \mult1_un159_sum_1_SUM[1] ), .D(\mult1_un159_sum_1_SUM[2] ), 
        .Y(un1_m8_1));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[14]  (.A(\i_s[14] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[14] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \un1_time1[7]  (.A(pulse_meash_0_tim[7]), 
        .B(\state[4]_net_1 ), .C(\mult1_un166_sum_1_SUM_RNIQ5884[1] ), 
        .Y(\un1_time1[7]_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_d  (.A(
        mult1_un201_sum_1_CO1), .B(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .C(
        \mult1_un194_sum_1_SUM[1] ), .Y(mult1_un201_sum_1_CO3_0_d));
    CFG3 #( .INIT(8'h69) )  \un24_k_v[0]  (.A(\valu[1]_net_1 ), .B(
        \mult1_un222_sum_1_SUM_0[4] ), .C(mult1_un222_sum_1_CO3), .Y(
        \un24_k_v[0]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_17[3]  (.A(
        un1_i_cry_22_S_0), .B(un1_i_cry_23_S_0), .C(un1_i_cry_24_S_0), 
        .D(un1_i_cry_25_S_0), .Y(\state_ns_i_a2_17[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \valu_RNO[12]  (.A(\state[4]_net_1 ), .B(
        pulse_meash_0_tim[12]), .Y(\valu_RNO[12]_net_1 ));
    SLE \valu[12]  (.D(\valu_RNO[12]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[12]_net_1 ));
    CFG3 #( .INIT(8'h06) )  \valu_RNI7VU53[5]  (.A(\valu[5]_net_1 ), 
        .B(mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .C(un1_N_5_i_2), .Y(
        un1_i3_mux_0));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_13 (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_12_net_1), .S(un1_i_cry_13_S_0), .Y(), .FCO(
        un1_i_cry_13_net_1));
    ARI1 #( .INIT(20'h65500) )  \i_cry[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[8]_net_1 ), .S(\i_s[9] ), .Y(), .FCO(\i_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[21]  (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[20]_net_1 ), .S(\i_s[21] ), .Y(), .FCO(
        \i_cry[21]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_bm[0]  (.A(\buff_2[0]_net_1 )
        , .B(\i[0]_net_1 ), .C(\buff_3[0]_net_1 ), .Y(
        \data_out_1_5_bm[0]_net_1 ));
    CFG4 #( .INIT(16'h3A30) )  \i_lm_0[0]  (.A(\i_cry_Y_0[0] ), .B(
        N_96), .C(\state[4]_net_1 ), .D(N_91), .Y(\i_lm[0] ));
    SLE \buff_3[1]  (.D(\k[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_3_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_3[1]_net_1 ));
    SLE \i[3]  (.D(\i_lm[3] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    CFG3 #( .INIT(8'h69) )  \valu_RNICB5V[13]  (.A(\valu[12]_net_1 ), 
        .B(un1_N_3_mux), .C(\valu[13]_net_1 ), .Y(
        \valu_RNICB5V[13]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[4]  (.A(\i_s[4] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[4] ));
    CFG3 #( .INIT(8'h45) )  \valu_RNI4LJS4[9]  (.A(\valu[9]_net_1 ), 
        .B(\valu[8]_net_1 ), .C(un1_N_5_1), .Y(mult1_un173_sum_1_CO1_0)
        );
    SLE \valu[2]  (.D(\un1_time1[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[2]_net_1 ));
    CFG4 #( .INIT(16'h7EBE) )  
        \un1_k_if_generate_plus.mult1_un194_sum_1_CO3_0_tz_0_1  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_1_RNO), .B(
        \mult1_un180_sum_1_SUM[4] ), .C(\valu[7]_net_1 ), .D(
        \mult1_un180_sum_1_SUM[2] ), .Y(mult1_un194_sum_1_CO3_0_tz_0_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_24 (.A(VCC_net_1), .B(
        \i[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_23_net_1), .S(un1_i_cry_24_S_0), .Y(), .FCO(
        un1_i_cry_24_net_1));
    CFG2 #( .INIT(4'h8) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_ANC2  (.A(
        mult1_un201_sum_1_CO1), .B(\mult1_un194_sum_1_SUM[1] ), .Y(
        mult1_un201_sum_1_ANC2));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_11 (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_10_net_1), .S(un1_i_cry_11_S_0), .Y(), .FCO(
        un1_i_cry_11_net_1));
    ARI1 #( .INIT(20'h65500) )  \i_cry[16]  (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[15]_net_1 ), .S(\i_s[16] ), .Y(), .FCO(
        \i_cry[16]_net_1 ));
    SLE \buff_5[4]  (.D(\k[5] ), .CLK(FCCC_0_GL0), .EN(
        buff_5_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\buff_5[5] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[7]_net_1 ), .S(\i_s[8] ), .Y(), .FCO(\i_cry[8]_net_1 ));
    CFG4 #( .INIT(16'h9024) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0_RNO_0  (.A(
        \valu[3]_net_1 ), .B(\valu[4]_net_1 ), .C(N_3560_i), .D(
        \mult1_un201_sum_1_SUM[4] ), .Y(mult1_un215_sum_1_ANC3_0_RNO_0)
        );
    ARI1 #( .INIT(20'h65500) )  \i_cry[0]  (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(GND_net_1), 
        .S(), .Y(\i_cry_Y_0[0] ), .FCO(\i_cry[0]_net_1 ));
    SLE \valu[1]  (.D(\un1_time1[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_i_a3_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \valu[1]_net_1 ));
    SLE \buff_2[4]  (.D(\k[5] ), .CLK(FCCC_0_GL0), .EN(
        buff_2_1_sqmuxa_1_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_2[5] ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_0_a2_14[5]  (.A(
        \i[7]_net_1 ), .B(\i[6]_net_1 ), .C(\i[4]_net_1 ), .D(
        \i[3]_net_1 ), .Y(\state_ns_i_0_a2_14[5]_net_1 ));
    CFG4 #( .INIT(16'hE44E) )  \un1_time1[3]  (.A(\state[4]_net_1 ), 
        .B(pulse_meash_0_tim[3]), .C(mult1_un201_sum_1_CO3), .D(
        \mult1_un201_sum_1_SUM_2[4] ), .Y(\un1_time1[3]_net_1 ));
    SLE \i[1]  (.D(\i_lm[1] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un173_sum_1_SUM[1]  (.A(
        \valu[9]_net_1 ), .B(\valu[8]_net_1 ), .C(
        mult1_un166_sum_1_CO3), .Y(\mult1_un173_sum_1_SUM[1] ));
    CFG4 #( .INIT(16'hDB24) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_tz_s_0_RNO_1  
        (.A(\valu[5]_net_1 ), .B(\valu[6]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[4] ), .D(\mult1_un187_sum_1_SUM[1] ), 
        .Y(d_N_19));
    CFG4 #( .INIT(16'h24DB) )  
        \un1_k_if_generate_plus.mult1_un166_sum_1_SUM[2]  (.A(
        \valu[9]_net_1 ), .B(\valu[10]_net_1 ), .C(
        \mult1_un159_sum_1_SUM[4] ), .D(\mult1_un159_sum_1_SUM[1] ), 
        .Y(\mult1_un166_sum_1_SUM[2] ));
    CFG2 #( .INIT(4'h4) )  \valu_RNIPTUG[4]  (.A(\valu[5]_net_1 ), .B(
        \valu[4]_net_1 ), .Y(d_m12_0_a3_0));
    CFG4 #( .INIT(16'h2000) )  \state_ns_i_a3_0[3]  (.A(N_90), .B(
        \state[1]_net_1 ), .C(\state_ns_i_a2[3]_net_1 ), .D(N_89), .Y(
        N_93));
    CFG4 #( .INIT(16'h05F3) )  \data_out_1_5_am_1_1[1]  (.A(
        \buff_1[1]_net_1 ), .B(\buff_0[1]_net_1 ), .C(\i[2]_net_1 ), 
        .D(\i[0]_net_1 ), .Y(\data_out_1_5_am_1_1[1]_net_1 ));
    CFG4 #( .INIT(16'hFAF8) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO3_0_0_1  (.A(
        mult1_un194_sum_1_CO3_0_tz_0_RNIU7S42), .B(
        mult1_un201_sum_1_CO2_0_d), .C(mult1_un201_sum_1_ANC3), .D(
        mult1_un201_sum_1_CO3_0_tz_s_0), .Y(
        mult1_un201_sum_1_CO3_0_0_1));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_0_a2_15[5]  (.A(
        \i[17]_net_1 ), .B(\i[16]_net_1 ), .C(\i[13]_net_1 ), .D(
        \i[12]_net_1 ), .Y(\state_ns_i_0_a2_15[5]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \state_ns_i_a2_13[3]  (.A(
        un1_i_cry_7_S_0), .B(un1_i_cry_8_S), .C(un1_i_cry_9_S_0), .D(
        un1_i_cry_10_S_0), .Y(\state_ns_i_a2_13[3]_net_1 ));
    SLE \buff_1[0]  (.D(\un1_angle[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        un1_rst_n_inv_2_i_0_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_1[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM_0[4]  (.A(
        \mult1_un215_sum_1_SUM_0_0[4] ), .B(un1_m6_1_0), .C(
        mult1_un208_sum_1_CO2), .D(un1_i2_mux), .Y(
        \mult1_un215_sum_1_SUM_0[4] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[22]  (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[21]_net_1 ), .S(\i_s[22] ), .Y(), .FCO(
        \i_cry[22]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[17]  (.A(\i_s[17] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[17] ));
    CFG3 #( .INIT(8'h1E) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_SUM[4]  (.A(
        mult1_un215_sum_1_CO3_0), .B(mult1_un215_sum_1_ANC3), .C(
        \mult1_un215_sum_1_SUM_0[4] ), .Y(\mult1_un215_sum_1_SUM[4] ));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[23]  (.A(\i_s[23] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[23] ));
    CFG3 #( .INIT(8'h69) )  
        \un1_k_if_generate_plus.mult1_un187_sum_1_SUM_0[4]  (.A(
        mult1_un180_sum_1_CO2), .B(\mult1_un180_sum_1_SUM_0[3] ), .C(
        \mult1_un180_sum_1_SUM[4] ), .Y(\mult1_un187_sum_1_SUM_0[4] ));
    ARI1 #( .INIT(20'h65500) )  \i_cry[19]  (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[18]_net_1 ), .S(\i_s[19] ), .Y(), .FCO(
        \i_cry[19]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_ns[2]  (.A(
        \data_out_1_5_am[2]_net_1 ), .B(\i[1]_net_1 ), .C(
        \data_out_1_5_bm[2]_net_1 ), .Y(\data_out_1[2] ));
    ARI1 #( .INIT(20'h4AA00) )  un1_i_cry_19 (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un1_i_cry_18_net_1), .S(un1_i_cry_19_S_0), .Y(), .FCO(
        un1_i_cry_19_net_1));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_bm[4]  (.A(\buff_2[5] ), .B(
        \i[0]_net_1 ), .C(\buff_3[5] ), .Y(\data_out_1_5_bm[4]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_1[0] ), .CLK(FCCC_0_GL0), .EN(
        data_out_0_sqmuxa), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        time_sender_0_data_out_0));
    SLE \i[18]  (.D(\i_lm[18] ), .CLK(FCCC_0_GL0), .EN(N_84_i_0), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[18]_net_1 ));
    CFG4 #( .INIT(16'h1428) )  \valu_RNI7QM15[7]  (.A(\valu[8]_net_1 ), 
        .B(\valu[7]_net_1 ), .C(\valu[6]_net_1 ), .D(
        \mult1_un166_sum_1_SUM_RNIQ5884[1] ), .Y(un1_i1_mux));
    CFG4 #( .INIT(16'hA030) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_CO3_0  (.A(
        \valu[2]_net_1 ), .B(mult1_un215_sum_1_CO3_0_RNO), .C(
        \mult1_un194_sum_1_SUM_RNIMGHHA[2] ), .D(un1_i5_mux_0), .Y(
        mult1_un215_sum_1_CO3_0));
    CFG2 #( .INIT(4'h2) )  \i_lm_0[15]  (.A(\i_s[15] ), .B(
        \un1_clk_inv_i_0_o3[0]_net_1 ), .Y(\i_lm[15] ));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un159_sum_1_SUM[1]  (.A(
        \valu[10]_net_1 ), .B(\valu_RNI32OE1[13]_net_1 ), .C(
        \valu[11]_net_1 ), .Y(\mult1_un159_sum_1_SUM[1] ));
    CFG3 #( .INIT(8'hE2) )  \data_out_1_5_ns[4]  (.A(
        \data_out_1_5_am[4]_net_1 ), .B(\i[1]_net_1 ), .C(
        \data_out_1_5_bm[4]_net_1 ), .Y(\data_out_1[5] ));
    CFG3 #( .INIT(8'hF6) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_CO1_1_RNO  (.A(
        \valu[4]_net_1 ), .B(\valu[5]_net_1 ), .C(
        \mult1_un187_sum_1_SUM[4] ), .Y(un1_m8_i_0));
    SLE \buff_5[2]  (.D(\k[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        buff_5_1_sqmuxa_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \buff_5[2]_net_1 ));
    CFG4 #( .INIT(16'h7DD7) )  
        \un1_k_if_generate_plus.mult1_un215_sum_1_ANC3_0_RNO_1  (.A(
        N_3560_i), .B(\mult1_un194_sum_1_SUM[2] ), .C(un1_m7_i_0_1), 
        .D(un1_N_8), .Y(un1_m7_i_0));
    CFG3 #( .INIT(8'h96) )  
        \un1_k_if_generate_plus.mult1_un201_sum_1_SUM_1_RNIS7JO[1]  (
        .A(\valu[3]_net_1 ), .B(\mult1_un201_sum_1_SUM_1[1] ), .C(
        mult1_un194_sum_1_ANC3_0_1), .Y(un1_N_5_i_2));
    
endmodule


module BT_module(
       BT_module_0_data_buf,
       rx_dout_reg,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       BT_module_0_oen,
       COREUART_0_RXRDY
    );
output [7:0] BT_module_0_data_buf;
input  [7:0] rx_dout_reg;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
output BT_module_0_oen;
input  COREUART_0_RXRDY;

    wire GND_net_1, \TX_RX_repiter[0]_net_1 , VCC_net_1, 
        \TX_RX_repiter_ns[0] , \TX_RX_repiter[1]_net_1 , N_19_i_0;
    
    SLE \data_buf[4]  (.D(rx_dout_reg[4]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[4]));
    SLE \TX_RX_repiter[1]  (.D(\TX_RX_repiter[0]_net_1 ), .CLK(
        FCCC_0_GL0), .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \TX_RX_repiter[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \data_buf[1]  (.D(rx_dout_reg[1]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[1]));
    SLE \data_buf[3]  (.D(rx_dout_reg[3]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[3]));
    CFG3 #( .INIT(8'h02) )  \TX_RX_repiter_ns_0_a2[0]  (.A(
        COREUART_0_RXRDY), .B(\TX_RX_repiter[1]_net_1 ), .C(
        \TX_RX_repiter[0]_net_1 ), .Y(\TX_RX_repiter_ns[0] ));
    SLE \data_buf[0]  (.D(rx_dout_reg[0]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[0]));
    VCC VCC (.Y(VCC_net_1));
    SLE \TX_RX_repiter[0]  (.D(\TX_RX_repiter_ns[0] ), .CLK(FCCC_0_GL0)
        , .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \TX_RX_repiter[0]_net_1 ));
    SLE \data_buf[6]  (.D(rx_dout_reg[6]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[6]));
    SLE \data_buf[5]  (.D(rx_dout_reg[5]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[5]));
    SLE oen (.D(\TX_RX_repiter[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        N_19_i_0), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(BT_module_0_oen));
    CFG2 #( .INIT(4'hE) )  oen_RNO (.A(\TX_RX_repiter[0]_net_1 ), .B(
        \TX_RX_repiter[1]_net_1 ), .Y(N_19_i_0));
    SLE \data_buf[7]  (.D(rx_dout_reg[7]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[7]));
    SLE \data_buf[2]  (.D(rx_dout_reg[2]), .CLK(FCCC_0_GL0), .EN(
        \TX_RX_repiter[0]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        BT_module_0_data_buf[2]));
    
endmodule


module servo_driver(
       FCCC_0_LOCK,
       FCCC_0_GL0,
       SERVO_PWM_c,
       un46_clk_0,
       un46_clk_1,
       un46_clk_2,
       un46_clk_3,
       N_234_0
    );
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
output SERVO_PWM_c;
input  un46_clk_0;
input  un46_clk_1;
input  un46_clk_2;
input  un46_clk_3;
input  N_234_0;

    wire un11_clk_13, VCC_net_1, un5_pulse_length_cry_12_S, 
        \state_d[2] , GND_net_1, un11_clk_14, 
        un5_pulse_length_cry_12_net_1, un11_clk_0, \P[0] , un11_clk_1, 
        un5_pulse_length_cry_0_Y, un11_clk_2, un5_pulse_length_cry_1_S, 
        un11_clk_3, un5_pulse_length_cry_2_S, un11_clk_4, 
        un5_pulse_length_cry_3_S, un11_clk_5, un5_pulse_length_cry_4_S, 
        un11_clk_6, un5_pulse_length_cry_5_S, un11_clk_7, 
        un5_pulse_length_cry_6_S, un11_clk_8, un5_pulse_length_cry_7_S, 
        un11_clk_9, un5_pulse_length_cry_8_S, un11_clk_10, 
        un5_pulse_length_cry_9_S, un11_clk_11, 
        un5_pulse_length_cry_10_S, un11_clk_12, 
        un5_pulse_length_cry_11_S, \state[0]_net_1 , N_67_i_0, 
        \state[1]_net_1 , \state_ns[1] , \state_d_i_0[2] , 
        \i[0]_net_1 , \i_lm[0] , \i[1]_net_1 , \i_lm[1] , \i[2]_net_1 , 
        \i_lm[2] , \i[3]_net_1 , \i_lm[3] , \i[4]_net_1 , \i_lm[4] , 
        \i[5]_net_1 , \i_lm[5] , \i[6]_net_1 , \i_lm[6] , \i[7]_net_1 , 
        \i_lm[7] , \i[8]_net_1 , \i_lm[8] , \i[9]_net_1 , \i_lm[9] , 
        \i[10]_net_1 , \i_lm[10] , \i[11]_net_1 , \i_lm[11] , 
        \i[12]_net_1 , \i_lm[12] , \i[13]_net_1 , \i_lm[13] , 
        \i[14]_net_1 , \i_lm[14] , \i[15]_net_1 , \i_lm[15] , 
        \i[16]_net_1 , \i_lm[16] , \i[17]_net_1 , \i_lm[17] , 
        \i[18]_net_1 , \i_lm[18] , \i[19]_net_1 , \i_lm[19] , 
        \i[20]_net_1 , \i_lm[20] , \i[21]_net_1 , \i_lm[21] , 
        \i[22]_net_1 , \i_lm[22] , \i[23]_net_1 , \i_lm[23] , 
        \i[24]_net_1 , \i_lm[24] , \i[25]_net_1 , \i_lm[25] , 
        \i[26]_net_1 , \i_lm[26] , \i[27]_net_1 , \i_lm[27] , 
        \i[28]_net_1 , \i_lm[28] , \i[29]_net_1 , \i_lm[29] , 
        \i[30]_net_1 , \i_lm[30] , un5_pulse_length_cry_0_net_1, 
        un5_pulse_length, un5_pulse_length_cry_1_net_1, \P[2] , 
        un5_pulse_length_cry_2_net_1, un5_pulse_length_axb_2, 
        un5_pulse_length_cry_3_net_1, un5_pulse_length_axb_3, 
        un5_pulse_length_cry_4_net_1, \P[5] , 
        un5_pulse_length_cry_5_net_1, un5_pulse_length_axb_5, 
        un5_pulse_length_cry_6_net_1, \P[7] , 
        un5_pulse_length_cry_7_net_1, un5_pulse_length_axb_7, 
        un5_pulse_length_cry_8_net_1, \P[9] , 
        un5_pulse_length_cry_9_net_1, \P[10] , 
        un5_pulse_length_cry_10_net_1, \P[11] , 
        un5_pulse_length_cry_11_net_1, un5_pulse_length_axb_11, 
        un5_pulse_length_axb_12, un11_clk_cry_3_net_1, 
        un11_clk_cry_4_net_1, un11_clk_cry_5_net_1, 
        un11_clk_cry_6_net_1, un11_clk_cry_7_net_1, 
        un11_clk_cry_8_net_1, un11_clk_cry_9_net_1, 
        un11_clk_cry_10_net_1, un11_clk_cry_11_net_1, 
        un11_clk_cry_12_net_1, un11_clk_cry_13_net_1, 
        un11_clk_cry_14_net_1, un11_clk_cry_15_net_1, 
        un11_clk_cry_16_net_1, un11_clk_cry_17_net_1, 
        un11_clk_cry_18_net_1, un11_clk_cry_19_net_1, 
        un11_clk_cry_20_net_1, un11_clk_cry_21_net_1, 
        un11_clk_cry_22_net_1, un11_clk_cry_23_net_1, 
        un11_clk_cry_24_net_1, un11_clk_cry_25_net_1, 
        un11_clk_cry_26_net_1, un11_clk_cry_27_net_1, 
        un11_clk_cry_28_net_1, un11_clk_cry_29_net_1, 
        un11_clk_cry_30_net_1, i_s_321_FCO, \i_cry[1]_net_1 , \i_s[1] , 
        \i_cry[2]_net_1 , \i_s[2] , \i_cry[3]_net_1 , \i_s[3] , 
        \i_cry[4]_net_1 , \i_s[4] , \i_cry[5]_net_1 , \i_s[5] , 
        \i_cry[6]_net_1 , \i_s[6] , \i_cry[7]_net_1 , \i_s[7] , 
        \i_cry[8]_net_1 , \i_s[8] , \i_cry[9]_net_1 , \i_s[9] , 
        \i_cry[10]_net_1 , \i_s[10] , \i_cry[11]_net_1 , \i_s[11] , 
        \i_cry[12]_net_1 , \i_s[12] , \i_cry[13]_net_1 , \i_s[13] , 
        \i_cry[14]_net_1 , \i_s[14] , \i_cry[15]_net_1 , \i_s[15] , 
        \i_cry[16]_net_1 , \i_s[16] , \i_cry[17]_net_1 , \i_s[17] , 
        \i_cry[18]_net_1 , \i_s[18] , \i_cry[19]_net_1 , \i_s[19] , 
        \i_cry[20]_net_1 , \i_s[20] , \i_cry[21]_net_1 , \i_s[21] , 
        \i_cry[22]_net_1 , \i_s[22] , \i_cry[23]_net_1 , \i_s[23] , 
        \i_cry[24]_net_1 , \i_s[24] , \i_cry[25]_net_1 , \i_s[25] , 
        \i_cry[26]_net_1 , \i_s[26] , \i_cry[27]_net_1 , \i_s[27] , 
        \i_cry[28]_net_1 , \i_s[28] , \i_s[30]_net_1 , 
        \i_cry[29]_net_1 , \i_s[29] , un1_state_0_sqmuxa_0_net_1, 
        un17_clklto30_7_net_1, un17_clklto30_6_net_1, 
        un17_clklto19_2_net_1, un17_clklto13_2_net_1, 
        un17_clklto30_8_net_1, un17_clklt13, un17_clklt19, 
        un17_clklto30_net_1;
    
    SLE \state[0]  (.D(N_67_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_4 (.A(VCC_net_1), 
        .B(\P[5] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_3_net_1), .S(un5_pulse_length_cry_4_S), 
        .Y(), .FCO(un5_pulse_length_cry_4_net_1));
    SLE \pulse_length[16]  (.D(un5_pulse_length_cry_12_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_13));
    SLE \i[7]  (.D(\i_lm[7] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    SLE \i[16]  (.D(\i_lm[16] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[16]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[14]  (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[13]_net_1 ), .S(\i_s[14] ), .Y(), .FCO(
        \i_cry[14]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_27 (.A(VCC_net_1), .B(
        \i[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_26_net_1), .S(), .Y(), .FCO(un11_clk_cry_27_net_1)
        );
    CFG2 #( .INIT(4'h8) )  \i_lm_0[24]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[24] ), .Y(\i_lm[24] ));
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_11 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_11), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un5_pulse_length_cry_10_net_1), .S(
        un5_pulse_length_cry_11_S), .Y(), .FCO(
        un5_pulse_length_cry_11_net_1));
    SLE \pulse_length[5]  (.D(un5_pulse_length_cry_1_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_2));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_20 (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_19_net_1), .S(), .Y(), .FCO(un11_clk_cry_20_net_1)
        );
    SLE \i[21]  (.D(\i_lm[21] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[21]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[20]  (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[19]_net_1 ), .S(\i_s[20] ), .Y(), .FCO(
        \i_cry[20]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_16 (.A(un11_clk_13), .B(
        \i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_15_net_1), .S(), .Y(), .FCO(un11_clk_cry_16_net_1)
        );
    SLE \i[0]  (.D(\i_lm[0] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    SLE \i[11]  (.D(\i_lm[11] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_13 (.A(un11_clk_10), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_12_net_1), .S(), .Y(), .FCO(un11_clk_cry_13_net_1)
        );
    CFG2 #( .INIT(4'h8) )  \i_lm_0[2]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[2] ), .Y(\i_lm[2] ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_24 (.A(VCC_net_1), .B(
        \i[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_23_net_1), .S(), .Y(), .FCO(un11_clk_cry_24_net_1)
        );
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_3 (.A(un11_clk_0), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(GND_net_1), 
        .S(), .Y(), .FCO(un11_clk_cry_3_net_1));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_18 (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_17_net_1), .S(), .Y(), .FCO(un11_clk_cry_18_net_1)
        );
    CFG4 #( .INIT(16'h5557) )  un17_clklto9 (.A(\i[9]_net_1 ), .B(
        \i[8]_net_1 ), .C(\i[7]_net_1 ), .D(\i[6]_net_1 ), .Y(
        un17_clklt13));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[27]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[27] ), .Y(\i_lm[27] ));
    CFG4 #( .INIT(16'h0001) )  un17_clklto30_7 (.A(\i[26]_net_1 ), .B(
        \i[25]_net_1 ), .C(\i[24]_net_1 ), .D(\i[23]_net_1 ), .Y(
        un17_clklto30_7_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[25]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[25] ), .Y(\i_lm[25] ));
    GND GND (.Y(GND_net_1));
    SLE \i[23]  (.D(\i_lm[23] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[23]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_12 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_12), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un5_pulse_length_cry_11_net_1), .S(
        un5_pulse_length_cry_12_S), .Y(), .FCO(
        un5_pulse_length_cry_12_net_1));
    CFG2 #( .INIT(4'h2) )  \i_RNO[0]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i[0]_net_1 ), .Y(\i_lm[0] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[23]  (.A(VCC_net_1), .B(
        \i[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[22]_net_1 ), .S(\i_s[23] ), .Y(), .FCO(
        \i_cry[23]_net_1 ));
    SLE \i[13]  (.D(\i_lm[13] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_7 (.A(un11_clk_4), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_6_net_1), .S(), .Y(), .FCO(un11_clk_cry_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[15]  (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[14]_net_1 ), .S(\i_s[15] ), .Y(), .FCO(
        \i_cry[15]_net_1 ));
    SLE \pulse_length[10]  (.D(un5_pulse_length_cry_6_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_7));
    SLE \i[27]  (.D(\i_lm[27] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[27]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_22 (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_21_net_1), .S(), .Y(), .FCO(un11_clk_cry_22_net_1)
        );
    SLE \pulse_length[14]  (.D(un5_pulse_length_cry_10_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_11));
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_2 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_2), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_1_net_1), .S(un5_pulse_length_cry_2_S), 
        .Y(), .FCO(un5_pulse_length_cry_2_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[10]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[10] ), .Y(\i_lm[10] ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_9 (.A(un11_clk_6), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_8_net_1), .S(), .Y(), .FCO(un11_clk_cry_9_net_1));
    SLE \i[17]  (.D(\i_lm[17] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[17]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un17_clklto13_2 (.A(\i[13]_net_1 ), .B(
        \i[12]_net_1 ), .C(\i[11]_net_1 ), .D(\i[10]_net_1 ), .Y(
        un17_clklto13_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[26]  (.A(VCC_net_1), .B(
        \i[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[25]_net_1 ), .S(\i_s[26] ), .Y(), .FCO(
        \i_cry[26]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[17]  (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[16]_net_1 ), .S(\i_s[17] ), .Y(), .FCO(
        \i_cry[17]_net_1 ));
    CFG4 #( .INIT(16'hA080) )  un17_clklto30 (.A(un17_clklto30_8_net_1)
        , .B(un17_clklt19), .C(un17_clklto30_7_net_1), .D(
        un17_clklto19_2_net_1), .Y(un17_clklto30_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[18]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[18] ), .Y(\i_lm[18] ));
    SLE \i[9]  (.D(\i_lm[9] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_0 (.A(VCC_net_1), 
        .B(un5_pulse_length), .C(GND_net_1), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(un5_pulse_length_cry_0_Y), .FCO(
        un5_pulse_length_cry_0_net_1));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_1 (.A(VCC_net_1), 
        .B(\P[2] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_0_net_1), .S(un5_pulse_length_cry_1_S), 
        .Y(), .FCO(un5_pulse_length_cry_1_net_1));
    SLE \pulse_length[8]  (.D(un5_pulse_length_cry_4_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_5));
    SLE \pulse_length[7]  (.D(un5_pulse_length_cry_3_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_4));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[29]  (.A(VCC_net_1), .B(
        \i[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[28]_net_1 ), .S(\i_s[29] ), .Y(), .FCO(
        \i_cry[29]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_26 (.A(VCC_net_1), .B(
        \i[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_25_net_1), .S(), .Y(), .FCO(un11_clk_cry_26_net_1)
        );
    SLE \pulse_length[13]  (.D(un5_pulse_length_cry_9_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_10));
    SLE \pulse_length[15]  (.D(un5_pulse_length_cry_11_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_12));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_19 (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_18_net_1), .S(), .Y(), .FCO(un11_clk_cry_19_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_5 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_5), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_4_net_1), .S(un5_pulse_length_cry_5_S), 
        .Y(), .FCO(un5_pulse_length_cry_5_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[11]  (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[10]_net_1 ), .S(\i_s[11] ), .Y(), .FCO(
        \i_cry[11]_net_1 ));
    SLE \i[25]  (.D(\i_lm[25] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[25]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_23 (.A(VCC_net_1), .B(
        \i[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_22_net_1), .S(), .Y(), .FCO(un11_clk_cry_23_net_1)
        );
    CFG4 #( .INIT(16'h0001) )  un17_clklto30_6 (.A(\i[30]_net_1 ), .B(
        \i[29]_net_1 ), .C(\i[28]_net_1 ), .D(\i[27]_net_1 ), .Y(
        un17_clklto30_6_net_1));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_8 (.A(VCC_net_1), 
        .B(\P[9] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_7_net_1), .S(un5_pulse_length_cry_8_S), 
        .Y(), .FCO(un5_pulse_length_cry_8_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[24]  (.A(VCC_net_1), .B(
        \i[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[23]_net_1 ), .S(\i_s[24] ), .Y(), .FCO(
        \i_cry[24]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[19]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[19] ), .Y(\i_lm[19] ));
    SLE \i[15]  (.D(\i_lm[15] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[15]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[3]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[3] ), .Y(\i_lm[3] ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[16]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[16] ), .Y(\i_lm[16] ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[20]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[20] ), .Y(\i_lm[20] ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_28 (.A(VCC_net_1), .B(
        \i[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_27_net_1), .S(), .Y(), .FCO(un11_clk_cry_28_net_1)
        );
    SLE \pulse_length[12]  (.D(un5_pulse_length_cry_8_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_9));
    MACC \un4_mulonly_0[31:18]  (.CLK({FCCC_0_GL0, FCCC_0_GL0}), .A({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, VCC_net_1, VCC_net_1, 
        GND_net_1, VCC_net_1, VCC_net_1, GND_net_1, VCC_net_1, 
        GND_net_1, VCC_net_1, VCC_net_1}), .A_EN({VCC_net_1, VCC_net_1})
        , .A_ARST_N({VCC_net_1, VCC_net_1}), .A_SRST_N({VCC_net_1, 
        VCC_net_1}), .B({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        un46_clk_3, un46_clk_2, un46_clk_1, un46_clk_0}), .B_EN({
        N_234_0, N_234_0}), .B_ARST_N({FCCC_0_LOCK, FCCC_0_LOCK}), 
        .B_SRST_N({VCC_net_1, VCC_net_1}), .C({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .C_EN({VCC_net_1, VCC_net_1}), 
        .C_ARST_N({VCC_net_1, VCC_net_1}), .C_SRST_N({VCC_net_1, 
        VCC_net_1}), .P_EN({VCC_net_1, VCC_net_1}), .P_ARST_N({
        VCC_net_1, VCC_net_1}), .P_SRST_N({VCC_net_1, VCC_net_1}), 
        .FDBKSEL(GND_net_1), .FDBKSEL_EN(VCC_net_1), .FDBKSEL_AL_N(
        VCC_net_1), .FDBKSEL_SL_N(VCC_net_1), .CDSEL(GND_net_1), 
        .CDSEL_EN(VCC_net_1), .CDSEL_AL_N(VCC_net_1), .CDSEL_SL_N(
        VCC_net_1), .ARSHFT17(GND_net_1), .ARSHFT17_EN(VCC_net_1), 
        .ARSHFT17_AL_N(VCC_net_1), .ARSHFT17_SL_N(VCC_net_1), .SUB(
        GND_net_1), .SUB_EN(VCC_net_1), .SUB_AL_N(VCC_net_1), 
        .SUB_SL_N(VCC_net_1), .CARRYIN(GND_net_1), .SIMD(GND_net_1), 
        .DOTP(GND_net_1), .OVFL_CARRYOUT_SEL(GND_net_1), .A_BYPASS({
        VCC_net_1, VCC_net_1}), .B_BYPASS({GND_net_1, GND_net_1}), 
        .C_BYPASS({VCC_net_1, VCC_net_1}), .P_BYPASS({VCC_net_1, 
        VCC_net_1}), .FDBKSEL_BYPASS(VCC_net_1), .FDBKSEL_AD(GND_net_1)
        , .FDBKSEL_SD_N(GND_net_1), .CDSEL_BYPASS(VCC_net_1), 
        .CDSEL_AD(GND_net_1), .CDSEL_SD_N(GND_net_1), .ARSHFT17_BYPASS(
        VCC_net_1), .ARSHFT17_AD(GND_net_1), .ARSHFT17_SD_N(GND_net_1), 
        .SUB_BYPASS(VCC_net_1), .SUB_AD(GND_net_1), .SUB_SD_N(
        GND_net_1), .CDIN({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .CDOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, 
        nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, nc19, nc20, 
        nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, 
        nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, nc39, nc40, 
        nc41, nc42, nc43}), .P({nc44, nc45, nc46, nc47, nc48, nc49, 
        nc50, nc51, nc52, nc53, nc54, nc55, nc56, nc57, nc58, nc59, 
        nc60, nc61, nc62, nc63, nc64, nc65, nc66, nc67, nc68, nc69, 
        nc70, nc71, nc72, nc73, un5_pulse_length_axb_12, 
        un5_pulse_length_axb_11, \P[11] , \P[10] , \P[9] , 
        un5_pulse_length_axb_7, \P[7] , un5_pulse_length_axb_5, \P[5] , 
        un5_pulse_length_axb_3, un5_pulse_length_axb_2, \P[2] , 
        un5_pulse_length, \P[0] }), .OVFL_CARRYOUT());
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_15 (.A(un11_clk_12), .B(
        \i[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_14_net_1), .S(), .Y(), .FCO(un11_clk_cry_15_net_1)
        );
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[6]_net_1 ), .S(\i_s[7] ), .Y(), .FCO(\i_cry[7]_net_1 ));
    SLE \i[22]  (.D(\i_lm[22] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[22]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_s[30]  (.A(VCC_net_1), .B(
        \i[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[29]_net_1 ), .S(\i_s[30]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[12]  (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[11]_net_1 ), .S(\i_s[12] ), .Y(), .FCO(
        \i_cry[12]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[6]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[6] ), .Y(\i_lm[6] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[18]  (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[17]_net_1 ), .S(\i_s[18] ), .Y(), .FCO(
        \i_cry[18]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  i_s_321 (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(i_s_321_FCO));
    SLE \i[2]  (.D(\i_lm[2] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    SLE \i[12]  (.D(\i_lm[12] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  un17_clklto30_8 (.A(\i[20]_net_1 ), .B(
        un17_clklto30_6_net_1), .C(\i[22]_net_1 ), .D(\i[21]_net_1 ), 
        .Y(un17_clklto30_8_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[28]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[28] ), .Y(\i_lm[28] ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_11 (.A(un11_clk_8), .B(
        \i[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_10_net_1), .S(), .Y(), .FCO(un11_clk_cry_11_net_1)
        );
    CFG2 #( .INIT(4'h8) )  \i_lm_0[1]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[1] ), .Y(\i_lm[1] ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[12]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[12] ), .Y(\i_lm[12] ));
    SLE \i[20]  (.D(\i_lm[20] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[20]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_9 (.A(VCC_net_1), 
        .B(\P[10] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_8_net_1), .S(un5_pulse_length_cry_9_S), 
        .Y(), .FCO(un5_pulse_length_cry_9_net_1));
    SLE \i[30]  (.D(\i_lm[30] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[30]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_6 (.A(VCC_net_1), 
        .B(\P[7] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_5_net_1), .S(un5_pulse_length_cry_6_S), 
        .Y(), .FCO(un5_pulse_length_cry_6_net_1));
    SLE \pulse_length[9]  (.D(un5_pulse_length_cry_5_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_6));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[11]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[11] ), .Y(\i_lm[11] ));
    SLE \i[10]  (.D(\i_lm[10] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    ARI1 #( .INIT(20'h65500) )  un5_pulse_length_cry_10 (.A(VCC_net_1), 
        .B(\P[11] ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_9_net_1), .S(un5_pulse_length_cry_10_S), 
        .Y(), .FCO(un5_pulse_length_cry_10_net_1));
    SLE \i[6]  (.D(\i_lm[6] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(i_s_321_FCO), 
        .S(\i_s[1] ), .Y(), .FCO(\i_cry[1]_net_1 ));
    SLE \i[29]  (.D(\i_lm[29] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[29]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[1]_net_1 ), .S(\i_s[2] ), .Y(), .FCO(\i_cry[2]_net_1 ));
    SLE \i[4]  (.D(\i_lm[4] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[10]  (.A(VCC_net_1), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[9]_net_1 ), .S(\i_s[10] ), .Y(), .FCO(\i_cry[10]_net_1 )
        );
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[5]_net_1 ), .S(\i_s[6] ), .Y(), .FCO(\i_cry[6]_net_1 ));
    SLE \pulse_length[6]  (.D(un5_pulse_length_cry_2_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_3));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[8]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[8] ), .Y(\i_lm[8] ));
    SLE \i[19]  (.D(\i_lm[19] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_3 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_3), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_2_net_1), .S(un5_pulse_length_cry_3_S), 
        .Y(), .FCO(un5_pulse_length_cry_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[25]  (.A(VCC_net_1), .B(
        \i[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[24]_net_1 ), .S(\i_s[25] ), .Y(), .FCO(
        \i_cry[25]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[29]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[29] ), .Y(\i_lm[29] ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_17 (.A(un11_clk_14), .B(
        \i[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_16_net_1), .S(), .Y(), .FCO(un11_clk_cry_17_net_1)
        );
    CFG2 #( .INIT(4'h8) )  \i_lm_0[26]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[26] ), .Y(\i_lm[26] ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_10 (.A(un11_clk_7), .B(
        \i[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_9_net_1), .S(), .Y(), .FCO(un11_clk_cry_10_net_1));
    SLE \i[24]  (.D(\i_lm[24] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[24]_net_1 ));
    CFG4 #( .INIT(16'h40EA) )  \state_ns_0[1]  (.A(\state[0]_net_1 ), 
        .B(\state[1]_net_1 ), .C(un17_clklto30_net_1), .D(
        un11_clk_cry_30_net_1), .Y(\state_ns[1] ));
    CFG4 #( .INIT(16'h5111) )  un17_clklto15 (.A(\i[15]_net_1 ), .B(
        \i[14]_net_1 ), .C(un17_clklto13_2_net_1), .D(un17_clklt13), 
        .Y(un17_clklt19));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[7]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[7] ), .Y(\i_lm[7] ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[13]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[13] ), .Y(\i_lm[13] ));
    SLE \i[14]  (.D(\i_lm[14] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[2]_net_1 ), .S(\i_s[3] ), .Y(), .FCO(\i_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[27]  (.A(VCC_net_1), .B(
        \i[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[26]_net_1 ), .S(\i_s[27] ), .Y(), .FCO(
        \i_cry[27]_net_1 ));
    SLE \pulse_length[4]  (.D(un5_pulse_length_cry_0_Y), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_1));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_29 (.A(VCC_net_1), .B(
        \i[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_28_net_1), .S(), .Y(), .FCO(un11_clk_cry_29_net_1)
        );
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_14 (.A(un11_clk_11), .B(
        \i[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_13_net_1), .S(), .Y(), .FCO(un11_clk_cry_14_net_1)
        );
    SLE \state[1]  (.D(\state_ns[1] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[30]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[30]_net_1 ), .Y(\i_lm[30] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[3]_net_1 ), .S(\i_s[4] ), .Y(), .FCO(\i_cry[4]_net_1 ));
    SLE \pulse_length[11]  (.D(un5_pulse_length_cry_7_S), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_8));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[22]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[22] ), .Y(\i_lm[22] ));
    SLE \i[5]  (.D(\i_lm[5] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_8 (.A(un11_clk_5), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_7_net_1), .S(), .Y(), .FCO(un11_clk_cry_8_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[9]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[9] ), .Y(\i_lm[9] ));
    SLE \i[8]  (.D(\i_lm[8] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    SLE \pulse_length[17]  (.D(un5_pulse_length_cry_12_net_1), .CLK(
        FCCC_0_GL0), .EN(\state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(un11_clk_14));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[21]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[21] ), .Y(\i_lm[21] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[13]  (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[12]_net_1 ), .S(\i_s[13] ), .Y(), .FCO(
        \i_cry[13]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[5]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[5] ), .Y(\i_lm[5] ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_5 (.A(un11_clk_2), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_4_net_1), .S(), .Y(), .FCO(un11_clk_cry_5_net_1));
    CFG3 #( .INIT(8'h0D) )  \state_RNO[0]  (.A(\state[0]_net_1 ), .B(
        un11_clk_cry_30_net_1), .C(\state[1]_net_1 ), .Y(N_67_i_0));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[14]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[14] ), .Y(\i_lm[14] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[4]_net_1 ), .S(\i_s[5] ), .Y(), .FCO(\i_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_6 (.A(un11_clk_3), .B(
        \i[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_5_net_1), .S(), .Y(), .FCO(un11_clk_cry_6_net_1));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_30 (.A(VCC_net_1), .B(
        \i[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_29_net_1), .S(), .Y(), .FCO(un11_clk_cry_30_net_1)
        );
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_25 (.A(VCC_net_1), .B(
        \i[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_24_net_1), .S(), .Y(), .FCO(un11_clk_cry_25_net_1)
        );
    CFG4 #( .INIT(16'h7FFF) )  un17_clklto19_2 (.A(\i[19]_net_1 ), .B(
        \i[18]_net_1 ), .C(\i[17]_net_1 ), .D(\i[16]_net_1 ), .Y(
        un17_clklto19_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[8]_net_1 ), .S(\i_s[9] ), .Y(), .FCO(\i_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[21]  (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[20]_net_1 ), .S(\i_s[21] ), .Y(), .FCO(
        \i_cry[21]_net_1 ));
    CFG2 #( .INIT(4'hE) )  state_s0_0_a3_i (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(\state_d_i_0[2] ));
    SLE \i[3]  (.D(\i_lm[3] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[4]  (.A(un1_state_0_sqmuxa_0_net_1), 
        .B(\i_s[4] ), .Y(\i_lm[4] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[16]  (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[15]_net_1 ), .S(\i_s[16] ), .Y(), .FCO(
        \i_cry[16]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[7]_net_1 ), .S(\i_s[8] ), .Y(), .FCO(\i_cry[8]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  un11_clk_cry_21 (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_20_net_1), .S(), .Y(), .FCO(un11_clk_cry_21_net_1)
        );
    SLE \pulse_length[3]  (.D(\P[0] ), .CLK(FCCC_0_GL0), .EN(
        \state_d[2] ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(un11_clk_0));
    SLE servo_pwm (.D(\state[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        \state_d_i_0[2] ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(SERVO_PWM_c));
    SLE \i[1]  (.D(\i_lm[1] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), .ALn(
        FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  un1_state_0_sqmuxa_0 (.A(
        \state[0]_net_1 ), .B(\state[1]_net_1 ), .C(
        un17_clklto30_net_1), .D(un11_clk_cry_30_net_1), .Y(
        un1_state_0_sqmuxa_0_net_1));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_12 (.A(un11_clk_9), .B(
        \i[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_11_net_1), .S(), .Y(), .FCO(un11_clk_cry_12_net_1)
        );
    SLE \i[28]  (.D(\i_lm[28] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[28]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un5_pulse_length_cry_7 (.A(VCC_net_1), 
        .B(un5_pulse_length_axb_7), .C(GND_net_1), .D(GND_net_1), .FCI(
        un5_pulse_length_cry_6_net_1), .S(un5_pulse_length_cry_7_S), 
        .Y(), .FCO(un5_pulse_length_cry_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[22]  (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[21]_net_1 ), .S(\i_s[22] ), .Y(), .FCO(
        \i_cry[22]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[17]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[17] ), .Y(\i_lm[17] ));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[23]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[23] ), .Y(\i_lm[23] ));
    CFG2 #( .INIT(4'h1) )  state_s0_0_a3 (.A(\state[0]_net_1 ), .B(
        \state[1]_net_1 ), .Y(\state_d[2] ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[19]  (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[18]_net_1 ), .S(\i_s[19] ), .Y(), .FCO(
        \i_cry[19]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \i_cry[28]  (.A(VCC_net_1), .B(
        \i[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \i_cry[27]_net_1 ), .S(\i_s[28] ), .Y(), .FCO(
        \i_cry[28]_net_1 ));
    SLE \i[18]  (.D(\i_lm[18] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[18]_net_1 ));
    ARI1 #( .INIT(20'h5AA55) )  un11_clk_cry_4 (.A(un11_clk_1), .B(
        \i[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un11_clk_cry_3_net_1), .S(), .Y(), .FCO(un11_clk_cry_4_net_1));
    CFG2 #( .INIT(4'h8) )  \i_lm_0[15]  (.A(un1_state_0_sqmuxa_0_net_1)
        , .B(\i_s[15] ), .Y(\i_lm[15] ));
    SLE \i[26]  (.D(\i_lm[26] ), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[26]_net_1 ));
    
endmodule


module Echo_control_COREUART_0_Rx_async_0s_1s_0s_1s_2s_3s(
       rx_byte,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       baud_clock,
       mss_sb_0_TX,
       stop_strobe,
       fifo_write,
       rx_idle
    );
output [7:0] rx_byte;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  baud_clock;
input  mss_sb_0_TX;
output stop_strobe;
output fifo_write;
output rx_idle;

    wire VCC_net_1, \rx_shift[3]_net_1 , rx_byte_1_sqmuxa, GND_net_1, 
        \rx_shift[4]_net_1 , \rx_shift[5]_net_1 , \rx_shift[6]_net_1 , 
        \rx_shift[7]_net_1 , \rx_bit_cnt[0]_net_1 , \rx_bit_cnt_4[0] , 
        \rx_bit_cnt[1]_net_1 , \rx_bit_cnt_4[1] , 
        \rx_bit_cnt[2]_net_1 , \rx_bit_cnt_4[2] , 
        \rx_bit_cnt[3]_net_1 , \rx_bit_cnt_4[3] , \rx_shift[1]_net_1 , 
        \rx_shift_11[1] , un1_samples7_1_0_net_1, \rx_shift[2]_net_1 , 
        \rx_shift_11[2] , \rx_shift_11[3] , \rx_shift_11[4] , 
        \rx_shift_11[5] , \rx_shift_11[6] , \rx_shift_11[7] , 
        \receive_count[0]_net_1 , N_182_i_0, \receive_count[1]_net_1 , 
        N_184_i_0, \receive_count[2]_net_1 , N_186_i_0, 
        \receive_count[3]_net_1 , N_188_i_0, \rx_shift[0]_net_1 , 
        \samples[0]_net_1 , \samples[1]_net_1 , \samples[2]_net_1 , 
        \rx_shift_11[0] , \rx_state[1]_net_1 , i9_mux_0, 
        \rx_statece[1]_net_1 , \rx_state[0]_net_1 , \rx_state_ns[0] , 
        framing_error_int_2_sqmuxa, \last_bit[0]_net_1 , 
        rx_state_0_sqmuxa, clear_parity_en_9_i_0, N_191, N_221, 
        rx_bit_cnt_0_sqmuxa, N_193, m16_am, m16_bm, rx_state19_NE_0, 
        clear_parity_en_9_3, \receive_count_3_i_a2_0_1[0] , N_24_mux, 
        N_22_mux, rx_state19_NE, rx_bit_cnt_1_sqmuxa, N_208, i5_mux, 
        CO1;
    
    CFG3 #( .INIT(8'h40) )  rx_bit_cnt_1_sqmuxa_0_a2 (.A(N_193), .B(
        \receive_count[3]_net_1 ), .C(baud_clock), .Y(
        rx_bit_cnt_1_sqmuxa));
    SLE \samples[0]  (.D(\samples[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[0]_net_1 ));
    SLE \rx_shift[2]  (.D(\rx_shift_11[2] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[2]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \rcv_cnt.receive_count_3_i_o2[0]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count_3_i_a2_0_1[0] ), .D(N_208), .Y(N_191));
    CFG3 #( .INIT(8'h08) )  \rcv_cnt.receive_count_3_i_a2_0_1_0[0]  (
        .A(\rx_state[1]_net_1 ), .B(\rx_state[0]_net_1 ), .C(
        \receive_count[3]_net_1 ), .Y(\receive_count_3_i_a2_0_1[0] ));
    CFG4 #( .INIT(16'h0200) )  rx_byte_1_sqmuxa_0_a2 (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .C(
        rx_state19_NE), .D(baud_clock), .Y(rx_byte_1_sqmuxa));
    CFG4 #( .INIT(16'hF0F8) )  un1_samples7_1_0 (.A(baud_clock), .B(
        \receive_count[3]_net_1 ), .C(rx_bit_cnt_0_sqmuxa), .D(N_193), 
        .Y(un1_samples7_1_0_net_1));
    SLE \rx_byte[0]  (.D(\rx_shift[0]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[0]));
    CFG4 #( .INIT(16'h0004) )  \rcv_cnt.receive_count_3_i_a2_0[3]  (.A(
        \receive_count[0]_net_1 ), .B(rx_idle), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_221));
    SLE \receive_count[1]  (.D(N_184_i_0), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[1]_net_1 ));
    CFG3 #( .INIT(8'hE4) )  \rx_state_ns_1_0_.m16_ns  (.A(
        \rx_state[1]_net_1 ), .B(m16_am), .C(m16_bm), .Y(
        \rx_state_ns[0] ));
    SLE \rx_shift[7]  (.D(\rx_shift_11[7] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[7]_net_1 ));
    CFG4 #( .INIT(16'hBFFF) )  fifo_write_RNO (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(
        clear_parity_en_9_3), .D(baud_clock), .Y(clear_parity_en_9_i_0)
        );
    SLE \rx_shift[0]  (.D(\rx_shift_11[0] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[0]  (.A(rx_idle), 
        .B(\rx_shift[1]_net_1 ), .Y(\rx_shift_11[0] ));
    SLE \receive_count[3]  (.D(N_188_i_0), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE fifo_write_inst_1 (.D(clear_parity_en_9_i_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(fifo_write));
    SLE \rx_byte[4]  (.D(\rx_shift[4]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[4]));
    CFG3 #( .INIT(8'hCA) )  \rx_state_ns_1_0_.m16_am  (.A(N_22_mux), 
        .B(rx_state19_NE), .C(\rx_state[0]_net_1 ), .Y(m16_am));
    SLE \rx_bit_cnt[2]  (.D(\rx_bit_cnt_4[2] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\rx_bit_cnt[2]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[3]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .C(CO1), .D(
        rx_bit_cnt_0_sqmuxa), .Y(\rx_bit_cnt_4[3] ));
    CFG2 #( .INIT(4'h8) )  rx_state_0_sqmuxa_0_a2 (.A(N_221), .B(
        \receive_count[3]_net_1 ), .Y(rx_state_0_sqmuxa));
    CFG3 #( .INIT(8'h04) )  rx_bit_cnt_0_sqmuxa_0_a2 (.A(
        \rx_state[0]_net_1 ), .B(baud_clock), .C(\rx_state[1]_net_1 ), 
        .Y(rx_bit_cnt_0_sqmuxa));
    SLE \rx_bit_cnt[1]  (.D(\rx_bit_cnt_4[1] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\rx_bit_cnt[1]_net_1 ));
    CFG2 #( .INIT(4'h1) )  rx_state_s0_0_a2 (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_idle));
    CFG4 #( .INIT(16'h0100) )  
        \receive_full_indicator.clear_parity_en_9_3  (.A(
        \rx_bit_cnt[1]_net_1 ), .B(\rx_bit_cnt[0]_net_1 ), .C(
        \rx_state[1]_net_1 ), .D(\rx_state[0]_net_1 ), .Y(
        clear_parity_en_9_3));
    CFG3 #( .INIT(8'h7F) )  \rcv_cnt.receive_count_3_i_o2[2]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .Y(N_193));
    CFG4 #( .INIT(16'h00E8) )  \receive_shift.rx_shift_11[7]  (.A(
        \samples[0]_net_1 ), .B(\samples[2]_net_1 ), .C(
        \samples[1]_net_1 ), .D(rx_idle), .Y(\rx_shift_11[7] ));
    CFG4 #( .INIT(16'h006A) )  \receive_count_RNO[2]  (.A(
        \receive_count[2]_net_1 ), .B(\receive_count[1]_net_1 ), .C(
        \receive_count[0]_net_1 ), .D(N_191), .Y(N_186_i_0));
    SLE stop_strobe_inst_1 (.D(framing_error_int_2_sqmuxa), .CLK(
        FCCC_0_GL0), .EN(baud_clock), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(stop_strobe));
    SLE \samples[1]  (.D(\samples[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[1]_net_1 ));
    CFG3 #( .INIT(8'hC5) )  \rx_state_ns_1_0_.m18  (.A(rx_state19_NE), 
        .B(i5_mux), .C(\rx_state[1]_net_1 ), .Y(i9_mux_0));
    SLE \rx_byte[1]  (.D(\rx_shift[1]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[1]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[2]  (.A(rx_idle), 
        .B(\rx_shift[3]_net_1 ), .Y(\rx_shift_11[2] ));
    SLE \receive_count[2]  (.D(N_186_i_0), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[2]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \un1_rx_bit_cnt_1.CO1  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_1_sqmuxa), .C(
        \rx_bit_cnt[1]_net_1 ), .Y(CO1));
    SLE \rx_state[1]  (.D(i9_mux_0), .CLK(FCCC_0_GL0), .EN(
        \rx_statece[1]_net_1 ), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[1]_net_1 ));
    SLE \rx_byte[6]  (.D(\rx_shift[6]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[6]));
    CFG3 #( .INIT(8'h06) )  \receive_count_RNO[1]  (.A(
        \receive_count[1]_net_1 ), .B(\receive_count[0]_net_1 ), .C(
        N_191), .Y(N_184_i_0));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h8) )  \rx_statece[1]  (.A(baud_clock), .B(
        \rx_state[0]_net_1 ), .Y(\rx_statece[1]_net_1 ));
    SLE \rx_shift[4]  (.D(\rx_shift_11[4] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[3]  (.A(rx_idle), 
        .B(\rx_shift[4]_net_1 ), .Y(\rx_shift_11[3] ));
    SLE \rx_byte[7]  (.D(\rx_shift[7]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[7]));
    CFG4 #( .INIT(16'hFFDE) )  \rcv_sm.rx_state19_NE  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_state19_NE_0), .C(
        \last_bit[0]_net_1 ), .D(\rx_bit_cnt[1]_net_1 ), .Y(
        rx_state19_NE));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[2]  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(CO1), .Y(
        \rx_bit_cnt_4[2] ));
    SLE \rx_byte[3]  (.D(\rx_shift[3]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[3]));
    CFG4 #( .INIT(16'h1000) )  \rx_state_ns_1_0_.m10  (.A(
        \receive_count[0]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_24_mux));
    CFG4 #( .INIT(16'h1001) )  \receive_count_RNO[3]  (.A(N_221), .B(
        N_208), .C(\receive_count[3]_net_1 ), .D(N_193), .Y(N_188_i_0));
    SLE \rx_byte[2]  (.D(\rx_shift[2]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[2]));
    CFG4 #( .INIT(16'h0103) )  \receive_count_RNO[0]  (.A(
        \receive_count[3]_net_1 ), .B(\receive_count[0]_net_1 ), .C(
        N_191), .D(N_221), .Y(N_182_i_0));
    SLE \rx_shift[6]  (.D(\rx_shift_11[6] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[6]_net_1 ));
    SLE \rx_shift[1]  (.D(\rx_shift_11[1] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[4]  (.A(rx_idle), 
        .B(\rx_shift[5]_net_1 ), .Y(\rx_shift_11[4] ));
    SLE \rx_shift[3]  (.D(\rx_shift_11[3] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[6]  (.A(rx_idle), 
        .B(\rx_shift[7]_net_1 ), .Y(\rx_shift_11[6] ));
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_state[0]_net_1 ));
    SLE \samples[2]  (.D(mss_sb_0_TX), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \samples[2]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  framing_error_int_2_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(\rx_state[0]_net_1 ), .C(
        \receive_count[3]_net_1 ), .D(N_193), .Y(
        framing_error_int_2_sqmuxa));
    SLE \receive_count[0]  (.D(N_182_i_0), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \receive_count[0]_net_1 ));
    SLE \rx_byte[5]  (.D(\rx_shift[5]_net_1 ), .CLK(FCCC_0_GL0), .EN(
        rx_byte_1_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_byte[5]));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[5]  (.A(rx_idle), 
        .B(\rx_shift[6]_net_1 ), .Y(\rx_shift_11[5] ));
    CFG4 #( .INIT(16'h0107) )  \rx_state_ns_1_0_.m14  (.A(
        \samples[2]_net_1 ), .B(\samples[0]_net_1 ), .C(N_24_mux), .D(
        \samples[1]_net_1 ), .Y(i5_mux));
    CFG3 #( .INIT(8'h12) )  \receive_shift.rx_bit_cnt_4[0]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(rx_bit_cnt_0_sqmuxa), .C(
        rx_bit_cnt_1_sqmuxa), .Y(\rx_bit_cnt_4[0] ));
    SLE \rx_shift[5]  (.D(\rx_shift_11[5] ), .CLK(FCCC_0_GL0), .EN(
        un1_samples7_1_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rx_shift[5]_net_1 ));
    CFG4 #( .INIT(16'hE800) )  \rcv_cnt.receive_count_3_i_a2[3]  (.A(
        \samples[0]_net_1 ), .B(\samples[2]_net_1 ), .C(
        \samples[1]_net_1 ), .D(rx_idle), .Y(N_208));
    SLE \rx_bit_cnt[0]  (.D(\rx_bit_cnt_4[0] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\rx_bit_cnt[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \receive_shift.rx_shift_11[1]  (.A(rx_idle), 
        .B(\rx_shift[2]_net_1 ), .Y(\rx_shift_11[1] ));
    CFG4 #( .INIT(16'h0004) )  \rx_state_ns_1_0_.m3  (.A(
        \receive_count[0]_net_1 ), .B(\receive_count[3]_net_1 ), .C(
        \receive_count[2]_net_1 ), .D(\receive_count[1]_net_1 ), .Y(
        N_22_mux));
    CFG4 #( .INIT(16'hC5C0) )  \rx_state_ns_1_0_.m16_bm  (.A(N_193), 
        .B(i5_mux), .C(\rx_state[0]_net_1 ), .D(
        \receive_count[3]_net_1 ), .Y(m16_bm));
    SLE \last_bit[0]  (.D(GND_net_1), .CLK(FCCC_0_GL0), .EN(
        rx_state_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \last_bit[0]_net_1 ));
    CFG2 #( .INIT(4'hB) )  \rcv_sm.rx_state19_NE_0  (.A(
        \rx_bit_cnt[2]_net_1 ), .B(\rx_bit_cnt[3]_net_1 ), .Y(
        rx_state19_NE_0));
    SLE \rx_bit_cnt[3]  (.D(\rx_bit_cnt_4[3] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\rx_bit_cnt[3]_net_1 ));
    CFG4 #( .INIT(16'h006C) )  \receive_shift.rx_bit_cnt_4[1]  (.A(
        \rx_bit_cnt[0]_net_1 ), .B(\rx_bit_cnt[1]_net_1 ), .C(
        rx_bit_cnt_1_sqmuxa), .D(rx_bit_cnt_0_sqmuxa), .Y(
        \rx_bit_cnt_4[1] ));
    
endmodule


module Echo_control_COREUART_0_ram128x8_pa4(
       data_out_0,
       rd_pointer,
       wr_pointer,
       tx_hold_reg_0,
       tx_hold_reg_1,
       tx_hold_reg_2,
       tx_hold_reg_3,
       tx_hold_reg_5,
       FCCC_0_GL0,
       fifo_write_tx
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  tx_hold_reg_0;
input  tx_hold_reg_1;
input  tx_hold_reg_2;
input  tx_hold_reg_3;
input  tx_hold_reg_5;
input  FCCC_0_GL0;
input  fifo_write_tx;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(FCCC_0_GL0), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(VCC_net_1), .A_DOUT_ARST_N(
        VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(VCC_net_1), 
        .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({rd_pointer[6], 
        rd_pointer[5], rd_pointer[4], rd_pointer[3], rd_pointer[2], 
        rd_pointer[1], rd_pointer[0], GND_net_1, GND_net_1, GND_net_1})
        , .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(VCC_net_1), 
        .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), 
        .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(VCC_net_1), 
        .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), .B_BLK({
        GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(FCCC_0_GL0), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        tx_hold_reg_5, tx_hold_reg_5, tx_hold_reg_3, tx_hold_reg_2, 
        tx_hold_reg_1, tx_hold_reg_0}), .C_WEN(INV_0_Y), .C_BLK({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_ADDR_LAT(
        GND_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .B_EN(GND_net_1), .B_ADDR_LAT(
        GND_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), .C_WIDTH({GND_net_1, 
        VCC_net_1, VCC_net_1}), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_tx), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module Echo_control_COREUART_0_fifo_ctrl_128_0s_128s_7s_8s(
       counter,
       tx_dout_reg,
       tx_hold_reg_0,
       tx_hold_reg_1,
       tx_hold_reg_2,
       tx_hold_reg_3,
       tx_hold_reg_5,
       fifo_write_tx,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_full_tx_i_0
    );
output [6:0] counter;
output [7:0] tx_dout_reg;
input  tx_hold_reg_0;
input  tx_hold_reg_1;
input  tx_hold_reg_2;
input  tx_hold_reg_3;
input  tx_hold_reg_5;
input  fifo_write_tx;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_full_tx_i_0;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , N_3820_i_0_net_1, 
        read_n_hold_net_1, read_n_hold_i_0, VCC_net_1, 
        un1_counter_cry_0_Y, GND_net_1, un1_counter_cry_1_0_S, 
        un1_counter_cry_2_0_S, un1_counter_cry_3_0_S, 
        un1_counter_cry_4_0_S, un1_counter_cry_5_0_S, 
        un1_counter_s_6_S, \data_out_0[4] , \data_out_0[5] , 
        \data_out_0[6] , \data_out_0[7] , \data_out_0[0] , 
        \data_out_0[1] , \data_out_0[2] , \data_out_0[3] , 
        \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_317_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_318_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        full_0_a2_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  full_0_a2_4_RNI02HF (.A(counter[0]), .B(
        full_0_a2_4_net_1), .C(counter[3]), .D(counter[2]), .Y(
        fifo_full_tx_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_318_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[2]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h5BB44) )  un1_counter_cry_2_0 (.A(counter[2]), 
        .B(fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        un1_counter_cry_1), .S(un1_counter_cry_2_0_S), .Y(), .FCO(
        un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[3])
        );
    SLE \counter[6]  (.D(un1_counter_s_6_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[6]));
    SLE read_n_hold (.D(fifo_read_tx), .CLK(FCCC_0_GL0), .EN(VCC_net_1)
        , .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h5BB44) )  un1_counter_cry_4_0 (.A(counter[4]), 
        .B(fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        un1_counter_cry_3), .S(un1_counter_cry_4_0_S), .Y(), .FCO(
        un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_317_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[7])
        );
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[4])
        );
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[4]));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[5]));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_318 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_318_FCO));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[5])
        );
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(FCCC_0_GL0), 
        .EN(N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[6]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  full_0_a2_4 (.A(counter[4]), .B(
        counter[5]), .C(counter[1]), .D(counter[6]), .Y(
        full_0_a2_4_net_1));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[0])
        );
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[1]));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[2])
        );
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[3]));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[6])
        );
    ARI1 #( .INIT(20'h5BB44) )  un1_counter_cry_3_0 (.A(counter[3]), 
        .B(fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        un1_counter_cry_2), .S(un1_counter_cry_3_0_S), .Y(), .FCO(
        un1_counter_cry_3));
    ARI1 #( .INIT(20'h59966) )  un1_counter_cry_0 (.A(counter[0]), .B(
        fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        GND_net_1), .S(), .Y(un1_counter_cry_0_Y), .FCO(
        un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(FCCC_0_GL0), .EN(
        N_3820_i_0_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(FCCC_0_GL0), 
        .EN(fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  N_3820_i_0 (.A(fifo_write_tx), .Y(
        N_3820_i_0_net_1));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNI6VUE (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    ARI1 #( .INIT(20'h5BB44) )  un1_counter_cry_1_0 (.A(counter[1]), 
        .B(fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        un1_counter_cry_0_net_1), .S(un1_counter_cry_1_0_S), .Y(), 
        .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(tx_dout_reg[1])
        );
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_317 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_317_FCO));
    ARI1 #( .INIT(20'h5BB44) )  un1_counter_cry_5_0 (.A(counter[5]), 
        .B(fifo_read_tx), .C(fifo_write_tx), .D(GND_net_1), .FCI(
        un1_counter_cry_4), .S(un1_counter_cry_5_0_S), .Y(), .FCO(
        un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_tx_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[4]_net_1 ));
    Echo_control_COREUART_0_ram128x8_pa4 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .tx_hold_reg_0(
        tx_hold_reg_0), .tx_hold_reg_1(tx_hold_reg_1), .tx_hold_reg_2(
        tx_hold_reg_2), .tx_hold_reg_3(tx_hold_reg_3), .tx_hold_reg_5(
        tx_hold_reg_5), .FCCC_0_GL0(FCCC_0_GL0), .fifo_write_tx(
        fifo_write_tx));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_tx_i_0), .C(fifo_write_tx), .D(counter[6]), .FCI(
        un1_counter_cry_5), .S(un1_counter_s_6_S), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter[0]));
    
endmodule


module Echo_control_COREUART_0_fifo_256x8_0s_4294967232s(
       counter,
       tx_dout_reg,
       tx_hold_reg_0,
       tx_hold_reg_1,
       tx_hold_reg_2,
       tx_hold_reg_3,
       tx_hold_reg_5,
       fifo_write_tx,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       fifo_read_tx,
       fifo_read_tx_i_0,
       fifo_full_tx_i_0
    );
output [6:0] counter;
output [7:0] tx_dout_reg;
input  tx_hold_reg_0;
input  tx_hold_reg_1;
input  tx_hold_reg_2;
input  tx_hold_reg_3;
input  tx_hold_reg_5;
input  fifo_write_tx;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  fifo_read_tx;
input  fifo_read_tx_i_0;
output fifo_full_tx_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    Echo_control_COREUART_0_fifo_ctrl_128_0s_128s_7s_8s 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.counter({counter[6], 
        counter[5], counter[4], counter[3], counter[2], counter[1], 
        counter[0]}), .tx_dout_reg({tx_dout_reg[7], tx_dout_reg[6], 
        tx_dout_reg[5], tx_dout_reg[4], tx_dout_reg[3], tx_dout_reg[2], 
        tx_dout_reg[1], tx_dout_reg[0]}), .tx_hold_reg_0(tx_hold_reg_0)
        , .tx_hold_reg_1(tx_hold_reg_1), .tx_hold_reg_2(tx_hold_reg_2), 
        .tx_hold_reg_3(tx_hold_reg_3), .tx_hold_reg_5(tx_hold_reg_5), 
        .fifo_write_tx(fifo_write_tx), .FCCC_0_LOCK(FCCC_0_LOCK), 
        .FCCC_0_GL0(FCCC_0_GL0), .fifo_read_tx(fifo_read_tx), 
        .fifo_read_tx_i_0(fifo_read_tx_i_0), .fifo_full_tx_i_0(
        fifo_full_tx_i_0));
    
endmodule


module Echo_control_COREUART_0_Tx_async_0s_1s_0s_1s_2s_3s_4s_5s_6s(
       tx_dout_reg,
       counter,
       fifo_read_tx,
       fifo_read_tx_i_0,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       xmit_pulse,
       Echo_control_0_TX,
       COREUART_0_TXRDY,
       fifo_full_tx_i_0,
       baud_clock,
       xmit_clock
    );
input  [7:0] tx_dout_reg;
input  [6:0] counter;
output fifo_read_tx;
output fifo_read_tx_i_0;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  xmit_pulse;
output Echo_control_0_TX;
output COREUART_0_TXRDY;
input  fifo_full_tx_i_0;
input  baud_clock;
input  xmit_clock;

    wire \tx_byte[2]_net_1 , VCC_net_1, N_119_i_0, GND_net_1, 
        \tx_byte[3]_net_1 , \tx_byte[4]_net_1 , \tx_byte[5]_net_1 , 
        \tx_byte[6]_net_1 , \tx_byte[7]_net_1 , 
        \xmit_bit_sel[0]_net_1 , \xmit_bit_sel_3[0] , 
        \xmit_bit_sel[1]_net_1 , N_111_i_0, \xmit_bit_sel[2]_net_1 , 
        N_113_i_0, \xmit_bit_sel[3]_net_1 , N_115_i_0, 
        \tx_byte[0]_net_1 , \tx_byte[1]_net_1 , tx_4_iv_i_a2, 
        N_129_i_0, fifo_read_en0_1_i_a3_i_net_1, \xmit_state[0]_net_1 , 
        \xmit_state_ns[0] , \xmit_state[1]_net_1 , 
        \xmit_state[6]_net_1 , \xmit_state[2]_net_1 , 
        \xmit_state_ns[2] , \xmit_state[3]_net_1 , N_101_i_0, 
        \xmit_state[5]_net_1 , \xmit_state_ns[5] , N_302_i_0, 
        \xmit_state_ns_0_a2_0_1[0]_net_1 , tx_2_u_i_m2_am_1_1, 
        tx_2_u_i_m2_am_1, tx_2_u_i_m2_bm_1_1, tx_2_u_i_m2_bm_1, 
        tx_2_u_i_m2_ns, N_328_3, N_326_5, \xmit_bit_sel_3_i_0_o2[3] , 
        \xmit_state_ns_0_a2[5]_net_1 ;
    
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_bm  (.A(
        \tx_byte[6]_net_1 ), .B(\tx_byte[7]_net_1 ), .C(
        tx_2_u_i_m2_bm_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_bm_1));
    SLE txrdy_int (.D(fifo_full_tx_i_0), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(COREUART_0_TXRDY));
    CFG3 #( .INIT(8'h7F) )  \xmit_cnt.xmit_bit_sel_3_i_0_o2[3]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[2]_net_1 ), .C(
        \xmit_bit_sel[0]_net_1 ), .Y(\xmit_bit_sel_3_i_0_o2[3] ));
    CFG3 #( .INIT(8'hE2) )  \xmit_sel.tx_2_u_i_m2_ns  (.A(
        tx_2_u_i_m2_am_1), .B(\xmit_bit_sel[2]_net_1 ), .C(
        tx_2_u_i_m2_bm_1), .Y(tx_2_u_i_m2_ns));
    SLE \xmit_state[3]  (.D(N_101_i_0), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_state[3]_net_1 ));
    SLE \tx_byte[0]  (.D(tx_dout_reg[0]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[0]_net_1 ));
    SLE \xmit_state[0]  (.D(\xmit_state_ns[0] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_state[0]_net_1 ));
    SLE \tx_byte[4]  (.D(tx_dout_reg[4]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \xmit_state_ns_0[5]  (.A(
        \xmit_state[5]_net_1 ), .B(xmit_pulse), .C(
        \xmit_state_ns_0_a2[5]_net_1 ), .Y(\xmit_state_ns[5] ));
    CFG3 #( .INIT(8'hAE) )  \xmit_state_ns_0[2]  (.A(
        \xmit_state[1]_net_1 ), .B(\xmit_state[2]_net_1 ), .C(
        xmit_pulse), .Y(\xmit_state_ns[2] ));
    CFG2 #( .INIT(4'h2) )  \xmit_cnt.xmit_bit_sel_3_a3_0_a2[0]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .Y(
        \xmit_bit_sel_3[0] ));
    CFG3 #( .INIT(8'h60) )  \xmit_bit_sel_RNO[1]  (.A(
        \xmit_bit_sel[1]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .Y(N_111_i_0));
    VCC VCC (.Y(VCC_net_1));
    SLE \tx_byte[5]  (.D(tx_dout_reg[5]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[5]_net_1 ));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_bm_1_1  (.A(
        \tx_byte[4]_net_1 ), .B(\tx_byte[5]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_bm_1_1));
    SLE \xmit_state[5]  (.D(\xmit_state_ns[5] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_state[5]_net_1 ));
    CFG3 #( .INIT(8'h51) )  \xmit_sel.tx_4_iv_i_a2  (.A(
        \xmit_state[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(
        tx_2_u_i_m2_ns), .Y(tx_4_iv_i_a2));
    CFG4 #( .INIT(16'h0020) )  \xmit_state_ns_0_a2[5]  (.A(
        \xmit_state[3]_net_1 ), .B(\xmit_bit_sel[3]_net_1 ), .C(
        xmit_pulse), .D(\xmit_bit_sel_3_i_0_o2[3] ), .Y(
        \xmit_state_ns_0_a2[5]_net_1 ));
    CFG4 #( .INIT(16'h8AAA) )  fifo_read_en0_1_i_a3_i_i (.A(
        \xmit_state[0]_net_1 ), .B(counter[5]), .C(N_328_3), .D(
        N_326_5), .Y(N_302_i_0));
    SLE \xmit_state[2]  (.D(\xmit_state_ns[2] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_state[2]_net_1 ));
    SLE \xmit_bit_sel[3]  (.D(N_115_i_0), .CLK(FCCC_0_GL0), .EN(
        xmit_pulse), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \xmit_state_RNIDBOR[2]  (.A(
        \xmit_state[2]_net_1 ), .B(baud_clock), .C(xmit_clock), .Y(
        N_119_i_0));
    CFG4 #( .INIT(16'hEAC0) )  \xmit_state_ns_0[0]  (.A(
        \xmit_state_ns_0_a2_0_1[0]_net_1 ), .B(\xmit_state[5]_net_1 ), 
        .C(xmit_pulse), .D(N_326_5), .Y(\xmit_state_ns[0] ));
    SLE \xmit_bit_sel[2]  (.D(N_113_i_0), .CLK(FCCC_0_GL0), .EN(
        xmit_pulse), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE tx (.D(tx_4_iv_i_a2), .CLK(FCCC_0_GL0), .EN(N_129_i_0), .ALn(
        FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(Echo_control_0_TX));
    SLE \tx_byte[3]  (.D(tx_dout_reg[3]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[3]_net_1 ));
    CFG4 #( .INIT(16'h0100) )  \xmit_state_ns_0_a2_0_1[0]  (.A(
        counter[6]), .B(counter[4]), .C(counter[5]), .D(
        \xmit_state[0]_net_1 ), .Y(\xmit_state_ns_0_a2_0_1[0]_net_1 ));
    SLE \tx_byte[7]  (.D(tx_dout_reg[7]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[7]_net_1 ));
    CFG4 #( .INIT(16'h00EC) )  \xmit_state_RNO[3]  (.A(
        \xmit_state[2]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(
        xmit_pulse), .D(\xmit_state_ns_0_a2[5]_net_1 ), .Y(N_101_i_0));
    CFG2 #( .INIT(4'h1) )  \xmit_state_ns_0_a2_0_3[0]  (.A(counter[4]), 
        .B(counter[6]), .Y(N_328_3));
    CFG4 #( .INIT(16'h60A0) )  \xmit_bit_sel_RNO[2]  (.A(
        \xmit_bit_sel[2]_net_1 ), .B(\xmit_bit_sel[0]_net_1 ), .C(
        \xmit_state[3]_net_1 ), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        N_113_i_0));
    CFG1 #( .INIT(2'h1) )  fifo_read_en0_RNIMOU (.A(fifo_read_tx), .Y(
        fifo_read_tx_i_0));
    SLE \tx_byte[6]  (.D(tx_dout_reg[6]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[6]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  fifo_read_en0_1_i_a3_i_a2_4 (.A(
        counter[3]), .B(counter[2]), .C(counter[1]), .D(counter[0]), 
        .Y(N_326_5));
    SLE \xmit_bit_sel[1]  (.D(N_111_i_0), .CLK(FCCC_0_GL0), .EN(
        xmit_pulse), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[1]_net_1 ));
    SLE \xmit_state[1]  (.D(\xmit_state[6]_net_1 ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_state[1]_net_1 ));
    SLE \xmit_bit_sel[0]  (.D(\xmit_bit_sel_3[0] ), .CLK(FCCC_0_GL0), 
        .EN(xmit_pulse), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \xmit_bit_sel[0]_net_1 ));
    SLE \tx_byte[2]  (.D(tx_dout_reg[2]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[2]_net_1 ));
    SLE fifo_read_en0 (.D(fifo_read_en0_1_i_a3_i_net_1), .CLK(
        FCCC_0_GL0), .EN(N_129_i_0), .ALn(FCCC_0_LOCK), .ADn(GND_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        fifo_read_tx));
    SLE \tx_byte[1]  (.D(tx_dout_reg[1]), .CLK(FCCC_0_GL0), .EN(
        N_119_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\tx_byte[1]_net_1 ));
    CFG3 #( .INIT(8'h84) )  \xmit_bit_sel_RNO[3]  (.A(
        \xmit_bit_sel[3]_net_1 ), .B(\xmit_state[3]_net_1 ), .C(
        \xmit_bit_sel_3_i_0_o2[3] ), .Y(N_115_i_0));
    CFG4 #( .INIT(16'h03F5) )  \xmit_sel.tx_2_u_i_m2_am_1_1  (.A(
        \tx_byte[0]_net_1 ), .B(\tx_byte[1]_net_1 ), .C(
        \xmit_bit_sel[1]_net_1 ), .D(\xmit_bit_sel[0]_net_1 ), .Y(
        tx_2_u_i_m2_am_1_1));
    SLE \xmit_state[6]  (.D(N_302_i_0), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_state[6]_net_1 ));
    CFG4 #( .INIT(16'h7555) )  fifo_read_en0_1_i_a3_i (.A(
        \xmit_state[0]_net_1 ), .B(counter[5]), .C(N_328_3), .D(
        N_326_5), .Y(fifo_read_en0_1_i_a3_i_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \xmit_state_RNIS58N1[1]  (.A(
        \xmit_state[0]_net_1 ), .B(\xmit_state[1]_net_1 ), .C(
        xmit_pulse), .D(\xmit_state[6]_net_1 ), .Y(N_129_i_0));
    CFG4 #( .INIT(16'hAC0F) )  \xmit_sel.tx_2_u_i_m2_am  (.A(
        \tx_byte[2]_net_1 ), .B(\tx_byte[3]_net_1 ), .C(
        tx_2_u_i_m2_am_1_1), .D(\xmit_bit_sel[1]_net_1 ), .Y(
        tx_2_u_i_m2_am_1));
    
endmodule


module Echo_control_COREUART_0_Clock_gen_0s_0s(
       xmit_clock,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       baud_clock,
       xmit_pulse
    );
output xmit_clock;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
output baud_clock;
output xmit_pulse;

    wire VCC_net_1, xmit_clock5, GND_net_1, \xmit_cntr[0]_net_1 , 
        \xmit_cntr_3[0] , \xmit_cntr[1]_net_1 , \xmit_cntr_3[1] , 
        \xmit_cntr[2]_net_1 , \xmit_cntr_3[2] , \xmit_cntr[3]_net_1 , 
        \xmit_cntr_3[3] , baud_cntr8_1_RNIEQ8C1_Y, \baud_cntr[0] , 
        \baud_cntr_s[0] , \baud_cntr[1] , \baud_cntr_s[1] , 
        \baud_cntr[2] , \baud_cntr_s[2] , \baud_cntr[3] , 
        \baud_cntr_s[3] , \baud_cntr[4] , \baud_cntr_s[4] , 
        \baud_cntr[5] , \baud_cntr_s[5] , \baud_cntr[6] , 
        \baud_cntr_s[6] , \baud_cntr[7] , \baud_cntr_s[7] , 
        \baud_cntr[8] , \baud_cntr_s[8] , \baud_cntr[9] , 
        \baud_cntr_s[9] , \baud_cntr[10] , \baud_cntr_s[10] , 
        \baud_cntr[11] , \baud_cntr_s[11] , \baud_cntr[12] , 
        \baud_cntr_s[12] , baud_cntr_cry_cy, baud_cntr8_8, 
        baud_cntr8_1, baud_cntr8_7, \baud_cntr_cry[0] , 
        \baud_cntr_cry[1] , \baud_cntr_cry[2] , \baud_cntr_cry[3] , 
        \baud_cntr_cry[4] , \baud_cntr_cry[5] , \baud_cntr_cry[6] , 
        \baud_cntr_cry[7] , \baud_cntr_cry[8] , \baud_cntr_cry[9] , 
        \baud_cntr_cry[10] , \baud_cntr_cry[11] , CO0;
    
    SLE \genblk1.baud_cntr[4]  (.D(\baud_cntr_s[4] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[4] )
        );
    SLE \genblk1.baud_cntr[1]  (.D(\baud_cntr_s[1] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[1] )
        );
    SLE \genblk1.baud_cntr[3]  (.D(\baud_cntr_s[3] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[3] )
        );
    SLE \xmit_cntr[3]  (.D(\xmit_cntr_3[3] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_cntr[3]_net_1 ));
    SLE \genblk1.baud_cntr[9]  (.D(\baud_cntr_s[9] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[9] )
        );
    SLE \genblk1.baud_clock_int  (.D(baud_cntr8_1_RNIEQ8C1_Y), .CLK(
        FCCC_0_GL0), .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        baud_clock));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_8  (
        .A(\baud_cntr[12] ), .B(\baud_cntr[7] ), .C(\baud_cntr[6] ), 
        .D(\baud_cntr[5] ), .Y(baud_cntr8_8));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI45C68[7]  (.A(
        VCC_net_1), .B(\baud_cntr[7] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[6] ), .S(\baud_cntr_s[7] ), .Y(), .FCO(
        \baud_cntr_cry[7] ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI3O1H7[5]  (.A(
        VCC_net_1), .B(\baud_cntr[5] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[4] ), .S(\baud_cntr_s[5] ), .Y(), .FCO(
        \baud_cntr_cry[5] ));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNIK6BB9[10]  (.A(
        VCC_net_1), .B(\baud_cntr[10] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[9] ), .S(\baud_cntr_s[10] ), .Y(), .FCO(
        \baud_cntr_cry[10] ));
    ARI1 #( .INIT(20'h44000) )  
        \genblk1.make_baud_cntr.baud_cntr8_1_RNIEQ8C1  (.A(
        baud_cntr8_8), .B(\baud_cntr[2] ), .C(baud_cntr8_1), .D(
        baud_cntr8_7), .FCI(VCC_net_1), .S(), .Y(
        baud_cntr8_1_RNIEQ8C1_Y), .FCO(baud_cntr_cry_cy));
    SLE \genblk1.baud_cntr[7]  (.D(\baud_cntr_s[7] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[7] )
        );
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI8QTM1[0]  (.A(
        VCC_net_1), .B(\baud_cntr[0] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(baud_cntr_cry_cy), .S(\baud_cntr_s[0] ), .Y(), .FCO(
        \baud_cntr_cry[0] ));
    SLE \genblk1.baud_cntr[5]  (.D(\baud_cntr_s[5] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[5] )
        );
    CFG4 #( .INIT(16'h8000) )  \make_xmit_clock.xmit_clock5  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[3]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(\xmit_cntr[0]_net_1 ), .Y(
        xmit_clock5));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6AAA) )  \make_xmit_clock.xmit_cntr_3_1.SUM[3]  
        (.A(\xmit_cntr[3]_net_1 ), .B(\xmit_cntr[2]_net_1 ), .C(
        \xmit_cntr[1]_net_1 ), .D(CO0), .Y(\xmit_cntr_3[3] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_1  (
        .A(\baud_cntr[4] ), .B(\baud_cntr[3] ), .C(\baud_cntr[1] ), .D(
        \baud_cntr[0] ), .Y(baud_cntr8_1));
    ARI1 #( .INIT(20'h61100) )  \genblk1.baud_cntr_RNI4JC67[4]  (.A(
        VCC_net_1), .B(baud_cntr8_1_RNIEQ8C1_Y), .C(\baud_cntr[4] ), 
        .D(GND_net_1), .FCI(\baud_cntr_cry[3] ), .S(\baud_cntr_s[4] ), 
        .Y(), .FCO(\baud_cntr_cry[4] ));
    SLE \genblk1.baud_cntr[8]  (.D(\baud_cntr_s[8] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[8] )
        );
    ARI1 #( .INIT(20'h61100) )  \genblk1.baud_cntr_RNIOKEF5[3]  (.A(
        VCC_net_1), .B(baud_cntr8_1_RNIEQ8C1_Y), .C(\baud_cntr[3] ), 
        .D(GND_net_1), .FCI(\baud_cntr_cry[2] ), .S(\baud_cntr_s[3] ), 
        .Y(), .FCO(\baud_cntr_cry[3] ));
    SLE \genblk1.baud_cntr[0]  (.D(\baud_cntr_s[0] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[0] )
        );
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI3UMR7[6]  (.A(
        VCC_net_1), .B(\baud_cntr[6] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[5] ), .S(\baud_cntr_s[6] ), .Y(), .FCO(
        \baud_cntr_cry[6] ));
    CFG4 #( .INIT(16'h0001) )  \genblk1.make_baud_cntr.baud_cntr8_7  (
        .A(\baud_cntr[11] ), .B(\baud_cntr[10] ), .C(\baud_cntr[9] ), 
        .D(\baud_cntr[8] ), .Y(baud_cntr8_7));
    ARI1 #( .INIT(20'h61100) )  \genblk1.baud_cntr_RNIHLRD3[1]  (.A(
        VCC_net_1), .B(baud_cntr8_1_RNIEQ8C1_Y), .C(\baud_cntr[1] ), 
        .D(GND_net_1), .FCI(\baud_cntr_cry[0] ), .S(\baud_cntr_s[1] ), 
        .Y(), .FCO(\baud_cntr_cry[1] ));
    SLE \xmit_cntr[2]  (.D(\xmit_cntr_3[2] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_cntr[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[1]  (.A(
        CO0), .B(\xmit_cntr[1]_net_1 ), .Y(\xmit_cntr_3[1] ));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI0OVQ9[11]  (.A(
        VCC_net_1), .B(\baud_cntr[11] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[10] ), .S(\baud_cntr_s[11] ), .Y(), .FCO(
        \baud_cntr_cry[11] ));
    SLE \genblk1.baud_cntr[10]  (.D(\baud_cntr_s[10] ), .CLK(
        FCCC_0_GL0), .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \baud_cntr[10] ));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNIDNGO3[2]  (.A(
        VCC_net_1), .B(\baud_cntr[2] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[1] ), .S(\baud_cntr_s[2] ), .Y(), .FCO(
        \baud_cntr_cry[2] ));
    SLE \genblk1.baud_cntr[6]  (.D(\baud_cntr_s[6] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[6] )
        );
    SLE xmit_clock_inst_1 (.D(xmit_clock5), .CLK(FCCC_0_GL0), .EN(
        baud_clock), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(xmit_clock));
    CFG2 #( .INIT(4'h8) )  \make_xmit_clock.xmit_cntr_3_1.CO0  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(CO0));
    ARI1 #( .INIT(20'h45500) )  \genblk1.baud_cntr_RNO[12]  (.A(
        VCC_net_1), .B(\baud_cntr[12] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[11] ), .S(\baud_cntr_s[12] ), .Y(), .FCO());
    SLE \genblk1.baud_cntr[12]  (.D(\baud_cntr_s[12] ), .CLK(
        FCCC_0_GL0), .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \baud_cntr[12] ));
    SLE \xmit_cntr[1]  (.D(\xmit_cntr_3[1] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_cntr[1]_net_1 ));
    SLE \genblk1.baud_cntr[2]  (.D(\baud_cntr_s[2] ), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\baud_cntr[2] )
        );
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI9MMR8[9]  (.A(
        VCC_net_1), .B(\baud_cntr[9] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[8] ), .S(\baud_cntr_s[9] ), .Y(), .FCO(
        \baud_cntr_cry[9] ));
    CFG2 #( .INIT(4'h8) )  xmit_pulse_inst_1 (.A(baud_clock), .B(
        xmit_clock), .Y(xmit_pulse));
    SLE \xmit_cntr[0]  (.D(\xmit_cntr_3[0] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\xmit_cntr[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \make_xmit_clock.xmit_cntr_3_1.SUM[0]  (.A(
        baud_clock), .B(\xmit_cntr[0]_net_1 ), .Y(\xmit_cntr_3[0] ));
    SLE \genblk1.baud_cntr[11]  (.D(\baud_cntr_s[11] ), .CLK(
        FCCC_0_GL0), .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \baud_cntr[11] ));
    CFG3 #( .INIT(8'h6A) )  \make_xmit_clock.xmit_cntr_3_1.SUM[2]  (.A(
        \xmit_cntr[2]_net_1 ), .B(\xmit_cntr[1]_net_1 ), .C(CO0), .Y(
        \xmit_cntr_3[2] ));
    ARI1 #( .INIT(20'h65500) )  \genblk1.baud_cntr_RNI6D1H8[8]  (.A(
        VCC_net_1), .B(\baud_cntr[8] ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\baud_cntr_cry[7] ), .S(\baud_cntr_s[8] ), .Y(), .FCO(
        \baud_cntr_cry[8] ));
    
endmodule


module Echo_control_COREUART_0_ram128x8_pa4_0(
       data_out_0,
       rd_pointer,
       wr_pointer,
       rx_byte,
       FCCC_0_GL0,
       fifo_write_rx_1
    );
output [7:0] data_out_0;
input  [6:0] rd_pointer;
input  [6:0] wr_pointer;
input  [7:0] rx_byte;
input  FCCC_0_GL0;
input  fifo_write_rx_1;

    wire VCC_net_1, GND_net_1, INV_0_Y;
    
    RAM64x18 RAM_128x8 (.A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, 
        nc7, nc8, nc9, data_out_0[7], data_out_0[6], data_out_0[5], 
        data_out_0[4], data_out_0[3], data_out_0[2], data_out_0[1], 
        data_out_0[0]}), .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27}), .BUSY(), .A_ADDR_CLK(FCCC_0_GL0), .A_DOUT_CLK(
        VCC_net_1), .A_ADDR_SRST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_ADDR_ARST_N(VCC_net_1), .A_DOUT_ARST_N(
        VCC_net_1), .A_ADDR_EN(VCC_net_1), .A_DOUT_EN(VCC_net_1), 
        .A_BLK({VCC_net_1, VCC_net_1}), .A_ADDR({rd_pointer[6], 
        rd_pointer[5], rd_pointer[4], rd_pointer[3], rd_pointer[2], 
        rd_pointer[1], rd_pointer[0], GND_net_1, GND_net_1, GND_net_1})
        , .B_ADDR_CLK(VCC_net_1), .B_DOUT_CLK(VCC_net_1), 
        .B_ADDR_SRST_N(VCC_net_1), .B_DOUT_SRST_N(VCC_net_1), 
        .B_ADDR_ARST_N(VCC_net_1), .B_DOUT_ARST_N(VCC_net_1), 
        .B_ADDR_EN(VCC_net_1), .B_DOUT_EN(VCC_net_1), .B_BLK({
        GND_net_1, GND_net_1}), .B_ADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .C_CLK(FCCC_0_GL0), .C_ADDR({
        wr_pointer[6], wr_pointer[5], wr_pointer[4], wr_pointer[3], 
        wr_pointer[2], wr_pointer[1], wr_pointer[0], GND_net_1, 
        GND_net_1, GND_net_1}), .C_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, rx_byte[7], rx_byte[6], 
        rx_byte[5], rx_byte[4], rx_byte[3], rx_byte[2], rx_byte[1], 
        rx_byte[0]}), .C_WEN(INV_0_Y), .C_BLK({VCC_net_1, VCC_net_1}), 
        .A_EN(VCC_net_1), .A_ADDR_LAT(GND_net_1), .A_DOUT_LAT(
        VCC_net_1), .A_WIDTH({GND_net_1, VCC_net_1, VCC_net_1}), .B_EN(
        GND_net_1), .B_ADDR_LAT(GND_net_1), .B_DOUT_LAT(VCC_net_1), 
        .B_WIDTH({GND_net_1, VCC_net_1, VCC_net_1}), .C_EN(VCC_net_1), 
        .C_WIDTH({GND_net_1, VCC_net_1, VCC_net_1}), .SII_LOCK(
        GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    INV INV_0 (.A(fifo_write_rx_1), .Y(INV_0_Y));
    GND GND (.Y(GND_net_1));
    
endmodule


module Echo_control_COREUART_0_fifo_ctrl_128_0s_128s_7s_8s_0(
       rx_dout,
       rx_byte,
       counter_0,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       N_3802_i_0,
       N_3803_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       full_0,
       full_4,
       fifo_empty_rx
    );
output [7:0] rx_dout;
input  [7:0] rx_byte;
output counter_0;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  N_3802_i_0;
input  N_3803_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output full_0;
output full_4;
output fifo_empty_rx;

    wire \rd_pointer[0]_net_1 , \rd_pointer_s[0] , 
        \wr_pointer[0]_net_1 , \wr_pointer_s[0] , read_n_hold_net_1, 
        read_n_hold_i_0, \counter[3]_net_1 , VCC_net_1, 
        un1_counter_cry_3_0_S_0, GND_net_1, \counter[4]_net_1 , 
        un1_counter_cry_4_0_S_0, \counter[5]_net_1 , 
        un1_counter_cry_5_0_S_0, \counter[6]_net_1 , 
        un1_counter_s_6_S_0, un1_counter_cry_0_Y_0, \counter[1]_net_1 , 
        un1_counter_cry_1_0_S_0, \counter[2]_net_1 , 
        un1_counter_cry_2_0_S_0, \data_out_0[0] , \data_out_0[1] , 
        \data_out_0[2] , \data_out_0[3] , \data_out_0[4] , 
        \data_out_0[5] , \data_out_0[6] , \data_out_0[7] , 
        \wr_pointer[1]_net_1 , \wr_pointer_s[1] , 
        \wr_pointer[2]_net_1 , \wr_pointer_s[2] , 
        \wr_pointer[3]_net_1 , \wr_pointer_s[3] , 
        \wr_pointer[4]_net_1 , \wr_pointer_s[4] , 
        \wr_pointer[5]_net_1 , \wr_pointer_s[5] , 
        \wr_pointer[6]_net_1 , \wr_pointer_s[6]_net_1 , 
        \rd_pointer[1]_net_1 , \rd_pointer_s[1] , 
        \rd_pointer[2]_net_1 , \rd_pointer_s[2] , 
        \rd_pointer[3]_net_1 , \rd_pointer_s[3] , 
        \rd_pointer[4]_net_1 , \rd_pointer_s[4] , 
        \rd_pointer[5]_net_1 , \rd_pointer_s[5] , 
        \rd_pointer[6]_net_1 , \rd_pointer_s[6]_net_1 , 
        un1_counter_cry_0_net_1, un1_counter_cry_1, un1_counter_cry_2, 
        un1_counter_cry_3, un1_counter_cry_4, un1_counter_cry_5, 
        rd_pointer_s_319_FCO, \rd_pointer_cry[1]_net_1 , 
        \rd_pointer_cry[2]_net_1 , \rd_pointer_cry[3]_net_1 , 
        \rd_pointer_cry[4]_net_1 , \rd_pointer_cry[5]_net_1 , 
        wr_pointer_s_320_FCO, \wr_pointer_cry[1]_net_1 , 
        \wr_pointer_cry[2]_net_1 , \wr_pointer_cry[3]_net_1 , 
        \wr_pointer_cry[4]_net_1 , \wr_pointer_cry[5]_net_1 , 
        empty_4_net_1;
    
    SLE \wr_pointer[5]  (.D(\wr_pointer_s[5] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  full_0_inst_1 (.A(\counter[1]_net_1 ), .B(
        \counter[2]_net_1 ), .Y(full_0));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[1]  (.A(VCC_net_1), .B(
        \wr_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        wr_pointer_s_320_FCO), .S(\wr_pointer_s[1] ), .Y(), .FCO(
        \wr_pointer_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[3]  (.A(VCC_net_1), .B(
        \wr_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[2]_net_1 ), .S(\wr_pointer_s[3] ), .Y(), .FCO(
        \wr_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[2]  (.A(VCC_net_1), .B(
        \wr_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[1]_net_1 ), .S(\wr_pointer_s[2] ), .Y(), .FCO(
        \wr_pointer_cry[2]_net_1 ));
    SLE \rd_pointer[2]  (.D(\rd_pointer_s[2] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[2]_net_1 ));
    SLE \counter[2]  (.D(un1_counter_cry_2_0_S_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[5]  (.A(VCC_net_1), .B(
        \wr_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[4]_net_1 ), .S(\wr_pointer_s[5] ), .Y(), .FCO(
        \wr_pointer_cry[5]_net_1 ));
    SLE \rd_pointer[5]  (.D(\rd_pointer_s[5] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[5]_net_1 ));
    ARI1 #( .INIT(20'h57788) )  un1_counter_cry_2_0 (.A(
        \counter[2]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(un1_counter_cry_1), .S(
        un1_counter_cry_2_0_S_0), .Y(), .FCO(un1_counter_cry_2));
    SLE \data_out[3]  (.D(\data_out_0[3] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[3]));
    SLE \counter[6]  (.D(un1_counter_s_6_S_0), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\counter[6]_net_1 ));
    SLE read_n_hold (.D(N_3802_i_0), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(read_n_hold_net_1));
    SLE \wr_pointer[1]  (.D(\wr_pointer_s[1] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_s[6]  (.A(VCC_net_1), .B(
        \rd_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[5]_net_1 ), .S(\rd_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h57788) )  un1_counter_cry_4_0 (.A(
        \counter[4]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(un1_counter_cry_3), .S(
        un1_counter_cry_4_0_S_0), .Y(), .FCO(un1_counter_cry_4));
    ARI1 #( .INIT(20'h4AA00) )  rd_pointer_s_319 (.A(VCC_net_1), .B(
        \rd_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(rd_pointer_s_319_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[1]  (.A(VCC_net_1), .B(
        \rd_pointer[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        rd_pointer_s_319_FCO), .S(\rd_pointer_s[1] ), .Y(), .FCO(
        \rd_pointer_cry[1]_net_1 ));
    SLE \data_out[7]  (.D(\data_out_0[7] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[7]));
    SLE \data_out[4]  (.D(\data_out_0[4] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[4]));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_s[6]  (.A(VCC_net_1), .B(
        \wr_pointer[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[5]_net_1 ), .S(\wr_pointer_s[6]_net_1 ), .Y(), 
        .FCO());
    SLE \wr_pointer[3]  (.D(\wr_pointer_s[3] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[3]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un1_counter_cry_4_0_S_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    SLE \counter[5]  (.D(un1_counter_cry_5_0_S_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    SLE \rd_pointer[0]  (.D(\rd_pointer_s[0] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[0]_net_1 ));
    SLE \data_out[5]  (.D(\data_out_0[5] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[5]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[3]  (.A(VCC_net_1), .B(
        \rd_pointer[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[2]_net_1 ), .S(\rd_pointer_s[3] ), .Y(), .FCO(
        \rd_pointer_cry[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  wr_pointer_s_320 (.A(VCC_net_1), .B(
        \wr_pointer[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(wr_pointer_s_320_FCO));
    ARI1 #( .INIT(20'h4AA00) )  \wr_pointer_cry[4]  (.A(VCC_net_1), .B(
        \wr_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \wr_pointer_cry[3]_net_1 ), .S(\wr_pointer_s[4] ), .Y(), .FCO(
        \wr_pointer_cry[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  \wr_pointer_RNO[0]  (.A(
        \wr_pointer[0]_net_1 ), .Y(\wr_pointer_s[0] ));
    SLE \wr_pointer[6]  (.D(\wr_pointer_s[6]_net_1 ), .CLK(FCCC_0_GL0), 
        .EN(N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[6]_net_1 ));
    SLE \data_out[0]  (.D(\data_out_0[0] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[0]));
    SLE \counter[1]  (.D(un1_counter_cry_1_0_S_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \wr_pointer[4]  (.D(\wr_pointer_s[4] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  read_n_hold_RNI58K5 (.A(read_n_hold_net_1), 
        .Y(read_n_hold_i_0));
    SLE \data_out[2]  (.D(\data_out_0[2] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[2]));
    SLE \counter[3]  (.D(un1_counter_cry_3_0_S_0), .CLK(FCCC_0_GL0), 
        .EN(VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \wr_pointer[0]  (.D(\wr_pointer_s[0] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[0]_net_1 ));
    SLE \data_out[6]  (.D(\data_out_0[6] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[6]));
    ARI1 #( .INIT(20'h57788) )  un1_counter_cry_3_0 (.A(
        \counter[3]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(un1_counter_cry_2), .S(
        un1_counter_cry_3_0_S_0), .Y(), .FCO(un1_counter_cry_3));
    ARI1 #( .INIT(20'h56699) )  un1_counter_cry_0 (.A(counter_0), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(GND_net_1), 
        .FCI(GND_net_1), .S(), .Y(un1_counter_cry_0_Y_0), .FCO(
        un1_counter_cry_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[5]  (.A(VCC_net_1), .B(
        \rd_pointer[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[4]_net_1 ), .S(\rd_pointer_s[5] ), .Y(), .FCO(
        \rd_pointer_cry[5]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  empty (.A(counter_0), .B(empty_4_net_1), 
        .C(\counter[2]_net_1 ), .D(\counter[1]_net_1 ), .Y(
        fifo_empty_rx));
    SLE \wr_pointer[2]  (.D(\wr_pointer_s[2] ), .CLK(FCCC_0_GL0), .EN(
        N_3803_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \wr_pointer[2]_net_1 ));
    SLE \rd_pointer[6]  (.D(\rd_pointer_s[6]_net_1 ), .CLK(FCCC_0_GL0), 
        .EN(fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[6]_net_1 ));
    SLE \rd_pointer[1]  (.D(\rd_pointer_s[1] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[1]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  empty_4 (.A(\counter[6]_net_1 ), .B(
        \counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(empty_4_net_1));
    ARI1 #( .INIT(20'h57788) )  un1_counter_cry_1_0 (.A(
        \counter[1]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(un1_counter_cry_0_net_1), 
        .S(un1_counter_cry_1_0_S_0), .Y(), .FCO(un1_counter_cry_1));
    CFG1 #( .INIT(2'h1) )  \rd_pointer_RNO[0]  (.A(
        \rd_pointer[0]_net_1 ), .Y(\rd_pointer_s[0] ));
    SLE \rd_pointer[3]  (.D(\rd_pointer_s[3] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[3]_net_1 ));
    SLE \data_out[1]  (.D(\data_out_0[1] ), .CLK(FCCC_0_GL0), .EN(
        read_n_hold_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout[1]));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[2]  (.A(VCC_net_1), .B(
        \rd_pointer[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[1]_net_1 ), .S(\rd_pointer_s[2] ), .Y(), .FCO(
        \rd_pointer_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h57788) )  un1_counter_cry_5_0 (.A(
        \counter[5]_net_1 ), .B(fifo_read_rx_0_sqmuxa), .C(
        fifo_write_rx_1), .D(GND_net_1), .FCI(un1_counter_cry_4), .S(
        un1_counter_cry_5_0_S_0), .Y(), .FCO(un1_counter_cry_5));
    SLE \rd_pointer[4]  (.D(\rd_pointer_s[4] ), .CLK(FCCC_0_GL0), .EN(
        fifo_read_rx_0_sqmuxa), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \rd_pointer[4]_net_1 ));
    Echo_control_COREUART_0_ram128x8_pa4_0 ram128_8_pa4 (.data_out_0({
        \data_out_0[7] , \data_out_0[6] , \data_out_0[5] , 
        \data_out_0[4] , \data_out_0[3] , \data_out_0[2] , 
        \data_out_0[1] , \data_out_0[0] }), .rd_pointer({
        \rd_pointer[6]_net_1 , \rd_pointer[5]_net_1 , 
        \rd_pointer[4]_net_1 , \rd_pointer[3]_net_1 , 
        \rd_pointer[2]_net_1 , \rd_pointer[1]_net_1 , 
        \rd_pointer[0]_net_1 }), .wr_pointer({\wr_pointer[6]_net_1 , 
        \wr_pointer[5]_net_1 , \wr_pointer[4]_net_1 , 
        \wr_pointer[3]_net_1 , \wr_pointer[2]_net_1 , 
        \wr_pointer[1]_net_1 , \wr_pointer[0]_net_1 }), .rx_byte({
        rx_byte[7], rx_byte[6], rx_byte[5], rx_byte[4], rx_byte[3], 
        rx_byte[2], rx_byte[1], rx_byte[0]}), .FCCC_0_GL0(FCCC_0_GL0), 
        .fifo_write_rx_1(fifo_write_rx_1));
    ARI1 #( .INIT(20'h4AA00) )  \rd_pointer_cry[4]  (.A(VCC_net_1), .B(
        \rd_pointer[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \rd_pointer_cry[3]_net_1 ), .S(\rd_pointer_s[4] ), .Y(), .FCO(
        \rd_pointer_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h47800) )  un1_counter_s_6 (.A(VCC_net_1), .B(
        fifo_read_rx_0_sqmuxa), .C(fifo_write_rx_1), .D(
        \counter[6]_net_1 ), .FCI(un1_counter_cry_5), .S(
        un1_counter_s_6_S_0), .Y(), .FCO());
    SLE \counter[0]  (.D(un1_counter_cry_0_Y_0), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(counter_0));
    CFG4 #( .INIT(16'h8000) )  full_4_inst_1 (.A(\counter[6]_net_1 ), 
        .B(\counter[5]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(full_4));
    
endmodule


module Echo_control_COREUART_0_fifo_256x8_0s_4294967232s_0(
       counter,
       rx_dout,
       rx_byte,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       N_3802_i_0,
       N_3803_i_0,
       fifo_read_rx_0_sqmuxa,
       fifo_write_rx_1,
       full_0,
       full_4,
       fifo_empty_rx
    );
output [0:0] counter;
output [7:0] rx_dout;
input  [7:0] rx_byte;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  N_3802_i_0;
input  N_3803_i_0;
input  fifo_read_rx_0_sqmuxa;
input  fifo_write_rx_1;
output full_0;
output full_4;
output fifo_empty_rx;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    Echo_control_COREUART_0_fifo_ctrl_128_0s_128s_7s_8s_0 
        CoreUART_top_COREUART_0_fifo_128x8_pa4 (.rx_dout({rx_dout[7], 
        rx_dout[6], rx_dout[5], rx_dout[4], rx_dout[3], rx_dout[2], 
        rx_dout[1], rx_dout[0]}), .rx_byte({rx_byte[7], rx_byte[6], 
        rx_byte[5], rx_byte[4], rx_byte[3], rx_byte[2], rx_byte[1], 
        rx_byte[0]}), .counter_0(counter[0]), .FCCC_0_LOCK(FCCC_0_LOCK)
        , .FCCC_0_GL0(FCCC_0_GL0), .N_3802_i_0(N_3802_i_0), 
        .N_3803_i_0(N_3803_i_0), .fifo_read_rx_0_sqmuxa(
        fifo_read_rx_0_sqmuxa), .fifo_write_rx_1(fifo_write_rx_1), 
        .full_0(full_0), .full_4(full_4), .fifo_empty_rx(fifo_empty_rx)
        );
    
endmodule


module Echo_control_COREUART_0_COREUART_1s_1s_0s_19s_0s_0s(
       rx_dout_reg,
       time_sender_0_data_out_0,
       time_sender_0_data_out_1,
       time_sender_0_data_out_2,
       time_sender_0_data_out_3,
       time_sender_0_data_out_5,
       FCCC_0_LOCK,
       FCCC_0_GL0,
       LED_3_c_i_0,
       COREUART_0_RXRDY,
       LED_3_c,
       BT_module_0_oen,
       Echo_control_0_TX,
       COREUART_0_TXRDY,
       mss_sb_0_TX
    );
output [7:0] rx_dout_reg;
input  time_sender_0_data_out_0;
input  time_sender_0_data_out_1;
input  time_sender_0_data_out_2;
input  time_sender_0_data_out_3;
input  time_sender_0_data_out_5;
input  FCCC_0_LOCK;
input  FCCC_0_GL0;
input  LED_3_c_i_0;
output COREUART_0_RXRDY;
input  LED_3_c;
input  BT_module_0_oen;
output Echo_control_0_TX;
output COREUART_0_TXRDY;
input  mss_sb_0_TX;

    wire rx_dout_reg_empty_net_1, rx_dout_reg_empty_i_0, VCC_net_1, 
        \rx_dout[5] , rx_dout_reg4_i_0, GND_net_1, \rx_dout[6] , 
        \rx_dout[7] , \tx_hold_reg[0]_net_1 , \tx_hold_reg[1]_net_1 , 
        \tx_hold_reg[2]_net_1 , \tx_hold_reg[3]_net_1 , 
        \tx_hold_reg[5] , \rx_dout[0] , \rx_dout[1] , \rx_dout[2] , 
        \rx_dout[3] , \rx_dout[4] , \rx_state[1]_net_1 , N_176_i, 
        rx_dout_reg4, rx_dout_reg_empty_1_sqmuxa_i_0, RXRDY5, 
        fifo_write_tx_net_1, \rx_state[0]_net_1 , \rx_state_ns[0] , 
        fifo_empty_rx, N_3802_i_0, fifo_write, \counter[0] , full_0, 
        full_4, N_3803_i_0, rx_idle, stop_strobe, 
        fifo_write_rx_1_net_1, fifo_read_rx_0_sqmuxa, xmit_clock, 
        baud_clock, xmit_pulse, \tx_dout_reg[0] , \tx_dout_reg[1] , 
        \tx_dout_reg[2] , \tx_dout_reg[3] , \tx_dout_reg[4] , 
        \tx_dout_reg[5] , \tx_dout_reg[6] , \tx_dout_reg[7] , 
        \counter_0[0] , \counter[1] , \counter[2] , \counter[3] , 
        \counter[4] , \counter[5] , \counter[6] , fifo_read_tx, 
        fifo_read_tx_i_0, fifo_full_tx_i_0, \rx_byte[0] , \rx_byte[1] , 
        \rx_byte[2] , \rx_byte[3] , \rx_byte[4] , \rx_byte[5] , 
        \rx_byte[6] , \rx_byte[7] ;
    
    CFG4 #( .INIT(16'h1555) )  fifo_write_rx_1_i (.A(fifo_write), .B(
        \counter[0] ), .C(full_0), .D(full_4), .Y(N_3803_i_0));
    SLE \rx_dout_reg[0]  (.D(\rx_dout[0] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[0])
        );
    CFG4 #( .INIT(16'hFFFB) )  fifo_read_rx_0_sqmuxa_0_a2_i (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(N_3802_i_0));
    CFG2 #( .INIT(4'h6) )  \rx_state_ns_0_x3[1]  (.A(
        \rx_state[0]_net_1 ), .B(\rx_state[1]_net_1 ), .Y(N_176_i));
    CFG4 #( .INIT(16'hEAAA) )  fifo_write_rx_1 (.A(fifo_write), .B(
        \counter[0] ), .C(full_0), .D(full_4), .Y(
        fifo_write_rx_1_net_1));
    Echo_control_COREUART_0_Rx_async_0s_1s_0s_1s_2s_3s make_RX (
        .rx_byte({\rx_byte[7] , \rx_byte[6] , \rx_byte[5] , 
        \rx_byte[4] , \rx_byte[3] , \rx_byte[2] , \rx_byte[1] , 
        \rx_byte[0] }), .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(
        FCCC_0_GL0), .baud_clock(baud_clock), .mss_sb_0_TX(mss_sb_0_TX)
        , .stop_strobe(stop_strobe), .fifo_write(fifo_write), .rx_idle(
        rx_idle));
    SLE \tx_hold_reg[0]  (.D(time_sender_0_data_out_0), .CLK(
        FCCC_0_GL0), .EN(LED_3_c_i_0), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\tx_hold_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h00AE) )  \rx_state_ns_0_a2[0]  (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(\rx_state_ns[0] ));
    SLE \rx_dout_reg[3]  (.D(\rx_dout[3] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[3])
        );
    Echo_control_COREUART_0_fifo_256x8_0s_4294967232s 
        \genblk2.tx_fifo  (.counter({\counter[6] , \counter[5] , 
        \counter[4] , \counter[3] , \counter[2] , \counter[1] , 
        \counter_0[0] }), .tx_dout_reg({\tx_dout_reg[7] , 
        \tx_dout_reg[6] , \tx_dout_reg[5] , \tx_dout_reg[4] , 
        \tx_dout_reg[3] , \tx_dout_reg[2] , \tx_dout_reg[1] , 
        \tx_dout_reg[0] }), .tx_hold_reg_0(\tx_hold_reg[0]_net_1 ), 
        .tx_hold_reg_1(\tx_hold_reg[1]_net_1 ), .tx_hold_reg_2(
        \tx_hold_reg[2]_net_1 ), .tx_hold_reg_3(\tx_hold_reg[3]_net_1 )
        , .tx_hold_reg_5(\tx_hold_reg[5] ), .fifo_write_tx(
        fifo_write_tx_net_1), .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(
        FCCC_0_GL0), .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .fifo_full_tx_i_0(fifo_full_tx_i_0));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg4_0 (.A(\rx_state[0]_net_1 ), .B(
        \rx_state[1]_net_1 ), .Y(rx_dout_reg4));
    SLE \tx_hold_reg[2]  (.D(time_sender_0_data_out_2), .CLK(
        FCCC_0_GL0), .EN(LED_3_c_i_0), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\tx_hold_reg[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  rx_dout_reg4_0_i (.A(\rx_state[0]_net_1 ), 
        .B(\rx_state[1]_net_1 ), .Y(rx_dout_reg4_i_0));
    SLE rx_dout_reg_empty (.D(rx_dout_reg4), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg_empty_1_sqmuxa_i_0), .ALn(FCCC_0_LOCK), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(rx_dout_reg_empty_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hFE) )  \genblk1.RXRDY5  (.A(rx_idle), .B(
        stop_strobe), .C(rx_dout_reg_empty_net_1), .Y(RXRDY5));
    CFG4 #( .INIT(16'h0004) )  fifo_read_rx_0_sqmuxa_0_a2 (.A(
        \rx_state[1]_net_1 ), .B(rx_dout_reg_empty_net_1), .C(
        fifo_empty_rx), .D(\rx_state[0]_net_1 ), .Y(
        fifo_read_rx_0_sqmuxa));
    Echo_control_COREUART_0_Tx_async_0s_1s_0s_1s_2s_3s_4s_5s_6s 
        make_TX (.tx_dout_reg({\tx_dout_reg[7] , \tx_dout_reg[6] , 
        \tx_dout_reg[5] , \tx_dout_reg[4] , \tx_dout_reg[3] , 
        \tx_dout_reg[2] , \tx_dout_reg[1] , \tx_dout_reg[0] }), 
        .counter({\counter[6] , \counter[5] , \counter[4] , 
        \counter[3] , \counter[2] , \counter[1] , \counter_0[0] }), 
        .fifo_read_tx(fifo_read_tx), .fifo_read_tx_i_0(
        fifo_read_tx_i_0), .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(
        FCCC_0_GL0), .xmit_pulse(xmit_pulse), .Echo_control_0_TX(
        Echo_control_0_TX), .COREUART_0_TXRDY(COREUART_0_TXRDY), 
        .fifo_full_tx_i_0(fifo_full_tx_i_0), .baud_clock(baud_clock), 
        .xmit_clock(xmit_clock));
    SLE \rx_dout_reg[4]  (.D(\rx_dout[4] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[4])
        );
    Echo_control_COREUART_0_Clock_gen_0s_0s make_CLOCK_GEN (
        .xmit_clock(xmit_clock), .FCCC_0_LOCK(FCCC_0_LOCK), 
        .FCCC_0_GL0(FCCC_0_GL0), .baud_clock(baud_clock), .xmit_pulse(
        xmit_pulse));
    SLE \rx_state[1]  (.D(N_176_i), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\rx_state[1]_net_1 ));
    SLE \rx_dout_reg[7]  (.D(\rx_dout[7] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[7])
        );
    GND GND (.Y(GND_net_1));
    SLE \rx_dout_reg[1]  (.D(\rx_dout[1] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[1])
        );
    SLE \rx_dout_reg[5]  (.D(\rx_dout[5] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[5])
        );
    CFG1 #( .INIT(2'h1) )  \genblk1.RXRDY_RNO  (.A(
        rx_dout_reg_empty_net_1), .Y(rx_dout_reg_empty_i_0));
    SLE \rx_dout_reg[6]  (.D(\rx_dout[6] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[6])
        );
    SLE \rx_state[0]  (.D(\rx_state_ns[0] ), .CLK(FCCC_0_GL0), .EN(
        VCC_net_1), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\rx_state[0]_net_1 ));
    SLE \genblk1.RXRDY  (.D(rx_dout_reg_empty_i_0), .CLK(FCCC_0_GL0), 
        .EN(RXRDY5), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        COREUART_0_RXRDY));
    Echo_control_COREUART_0_fifo_256x8_0s_4294967232s_0 
        \genblk3.rx_fifo  (.counter({\counter[0] }), .rx_dout({
        \rx_dout[7] , \rx_dout[6] , \rx_dout[5] , \rx_dout[4] , 
        \rx_dout[3] , \rx_dout[2] , \rx_dout[1] , \rx_dout[0] }), 
        .rx_byte({\rx_byte[7] , \rx_byte[6] , \rx_byte[5] , 
        \rx_byte[4] , \rx_byte[3] , \rx_byte[2] , \rx_byte[1] , 
        \rx_byte[0] }), .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(
        FCCC_0_GL0), .N_3802_i_0(N_3802_i_0), .N_3803_i_0(N_3803_i_0), 
        .fifo_read_rx_0_sqmuxa(fifo_read_rx_0_sqmuxa), 
        .fifo_write_rx_1(fifo_write_rx_1_net_1), .full_0(full_0), 
        .full_4(full_4), .fifo_empty_rx(fifo_empty_rx));
    SLE \tx_hold_reg[3]  (.D(time_sender_0_data_out_3), .CLK(
        FCCC_0_GL0), .EN(LED_3_c_i_0), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\tx_hold_reg[3]_net_1 ));
    SLE fifo_write_tx (.D(LED_3_c), .CLK(FCCC_0_GL0), .EN(VCC_net_1), 
        .ALn(FCCC_0_LOCK), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(fifo_write_tx_net_1));
    SLE \tx_hold_reg[1]  (.D(time_sender_0_data_out_1), .CLK(
        FCCC_0_GL0), .EN(LED_3_c_i_0), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\tx_hold_reg[1]_net_1 ));
    CFG2 #( .INIT(4'h7) )  rx_dout_reg_empty_1_sqmuxa_i (.A(
        rx_dout_reg4), .B(BT_module_0_oen), .Y(
        rx_dout_reg_empty_1_sqmuxa_i_0));
    SLE \rx_dout_reg[2]  (.D(\rx_dout[2] ), .CLK(FCCC_0_GL0), .EN(
        rx_dout_reg4_i_0), .ALn(FCCC_0_LOCK), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(rx_dout_reg[2])
        );
    SLE \tx_hold_reg[4]  (.D(time_sender_0_data_out_5), .CLK(
        FCCC_0_GL0), .EN(LED_3_c_i_0), .ALn(FCCC_0_LOCK), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\tx_hold_reg[5] ));
    
endmodule


module Echo_control_FCCC_0_FCCC(
       FCCC_0_LOCK,
       FCCC_0_GL0,
       OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC
    );
output FCCC_0_LOCK;
output FCCC_0_GL0;
input  OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC;

    wire LOCK, GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST (.A(GL0_net), .Y(FCCC_0_GL0));
    CCC #( .INIT(210'h0000007F88000045164000318C6318C1F18C61E80404040403100)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(LOCK), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(GND_net_1), .RCOSC_1MHZ(
        OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC), .XTLOSC(GND_net_1));
    CLKINT CCC_INST_RNIE1Q1 (.A(LOCK), .Y(FCCC_0_LOCK));
    
endmodule


module Echo_control_OSC_0_OSC(
       OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC
    );
output OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    RCOSC_1MHZ I_RCOSC_1MHZ (.CLKOUT(
        OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC));
    
endmodule


module delayer(
       FCCC_0_GL0,
       FCCC_0_LOCK,
       LED_2_c,
       pulse_meash_0_new_ready
    );
input  FCCC_0_GL0;
input  FCCC_0_LOCK;
output LED_2_c;
input  pulse_meash_0_new_ready;

    wire \i[16]_net_1 , VCC_net_1, \i_4[16] , GND_net_1, \i[17]_net_1 , 
        \i_4[17] , \i[18]_net_1 , \i_4[18] , \i[19]_net_1 , \i_4[19] , 
        \i[20]_net_1 , \i_4[20] , \i[21]_net_1 , \i_4[21] , 
        \i[22]_net_1 , \i_4[22] , \i[1]_net_1 , \i_4[1] , \i[2]_net_1 , 
        \i_4[2] , \i[3]_net_1 , \i_4[3] , \i[4]_net_1 , \i_4[4] , 
        \i[5]_net_1 , \i_4[5] , \i[6]_net_1 , \i_4[6] , \i[7]_net_1 , 
        \i_4[7] , \i[8]_net_1 , \i_4[8] , \i[9]_net_1 , \i_4[9] , 
        \i[10]_net_1 , \i_4[10] , \i[11]_net_1 , \i_4[11] , 
        \i[12]_net_1 , \i_4[12] , \i[13]_net_1 , \i_4[13] , 
        \i[14]_net_1 , \i_4[14] , \i[15]_net_1 , \i_4[15] , 
        \i[0]_net_1 , \i_4[0] , un9_clklto22_i_0_a3_RNI2GHT_Y, 
        i_4_cry_0_cy, un9_clklto22_i_0_a3_net_1, 
        un9_clklto22_i_0_a3_0_net_1, i_4_cry_0, i_4_cry_1, i_4_cry_2, 
        i_4_cry_3, i_4_cry_4, i_4_cry_5, i_4_cry_6, i_4_cry_7, 
        i_4_cry_8, i_4_cry_9, i_4_cry_10, i_4_cry_11, i_4_cry_12, 
        i_4_cry_13, i_4_cry_14, i_4_cry_15, i_4_cry_16, i_4_cry_17, 
        i_4_cry_18, i_4_cry_19, i_4_cry_20, i_4_cry_21, 
        un9_clklto22_i_0_a3_1_net_1, un9_clklto22_i_0_a2_2_3_net_1, 
        N_122, N_123, N_124, un9_clklto22_i_0_o2_net_1;
    
    ARI1 #( .INIT(20'h42200) )  \i_RNI64HF3[7]  (.A(VCC_net_1), .B(
        \i[7]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_6), .S(\i_4[7] ), .Y(), .FCO(i_4_cry_7));
    ARI1 #( .INIT(20'h42200) )  \i_RNIVAP71[0]  (.A(VCC_net_1), .B(
        \i[0]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_0_cy), .S(\i_4[0] ), .Y(), .FCO(i_4_cry_0));
    SLE \i[17]  (.D(\i_4[17] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[17]_net_1 ));
    CFG3 #( .INIT(8'h75) )  un9_clklto22_i_0_o2_0 (.A(\i[11]_net_1 ), 
        .B(\i[10]_net_1 ), .C(N_123), .Y(N_124));
    ARI1 #( .INIT(20'h42200) )  \i_RNIEFJ64[11]  (.A(VCC_net_1), .B(
        \i[11]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_10), .S(\i_4[11] ), .Y(), .FCO(i_4_cry_11));
    ARI1 #( .INIT(20'h4FFEF) )  un9_clklto22_i_0_a3_RNI2GHT (.A(
        pulse_meash_0_new_ready), .B(un9_clklto22_i_0_a3_net_1), .C(
        un9_clklto22_i_0_a3_0_net_1), .D(\i[22]_net_1 ), .FCI(
        VCC_net_1), .S(), .Y(un9_clklto22_i_0_a3_RNI2GHT_Y), .FCO(
        i_4_cry_0_cy));
    CFG3 #( .INIT(8'h01) )  un9_clklto22_i_0_a3_1 (.A(\i[17]_net_1 ), 
        .B(\i[16]_net_1 ), .C(\i[15]_net_1 ), .Y(
        un9_clklto22_i_0_a3_1_net_1));
    ARI1 #( .INIT(20'h42200) )  \i_RNI22953[6]  (.A(VCC_net_1), .B(
        \i[6]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_5), .S(\i_4[6] ), .Y(), .FCO(i_4_cry_6));
    SLE \i[21]  (.D(\i_4[21] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[21]_net_1 ));
    SLE \i[9]  (.D(\i_4[9] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[9]_net_1 ));
    SLE \i[2]  (.D(\i_4[2] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[2]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNO[22]  (.A(VCC_net_1), .B(
        \i[22]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_21), .S(\i_4[22] ), .Y(), .FCO());
    SLE \i[10]  (.D(\i_4[10] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[10]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIFN594[13]  (.A(VCC_net_1), .B(
        \i[13]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_12), .S(\i_4[13] ), .Y(), .FCO(i_4_cry_13));
    SLE \i[3]  (.D(\i_4[3] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[3]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNITJAE4[17]  (.A(VCC_net_1), .B(
        \i[17]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_16), .S(\i_4[17] ), .Y(), .FCO(i_4_cry_17));
    SLE \i[8]  (.D(\i_4[8] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[8]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIT61I1[1]  (.A(VCC_net_1), .B(
        \i[1]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_0), .S(\i_4[1] ), .Y(), .FCO(i_4_cry_1));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h42200) )  \i_RNI8B1D4[16]  (.A(VCC_net_1), .B(
        \i[16]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_15), .S(\i_4[16] ), .Y(), .FCO(i_4_cry_16));
    SLE \i[20]  (.D(\i_4[20] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[20]_net_1 ));
    SLE led (.D(un9_clklto22_i_0_a3_RNI2GHT_Y), .CLK(FCCC_0_GL0), .EN(
        FCCC_0_LOCK), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(LED_2_c));
    ARI1 #( .INIT(20'h42200) )  \i_RNIS39S1[2]  (.A(VCC_net_1), .B(
        \i[2]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_1), .S(\i_4[2] ), .Y(), .FCO(i_4_cry_2));
    ARI1 #( .INIT(20'h42200) )  \i_RNIUIS74[12]  (.A(VCC_net_1), .B(
        \i[12]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_11), .S(\i_4[12] ), .Y(), .FCO(i_4_cry_12));
    ARI1 #( .INIT(20'h42200) )  \i_RNIHB144[9]  (.A(VCC_net_1), .B(
        \i[9]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_8), .S(\i_4[9] ), .Y(), .FCO(i_4_cry_9));
    SLE \i[18]  (.D(\i_4[18] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[18]_net_1 ));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h42200) )  \i_RNIPB7I4[20]  (.A(VCC_net_1), .B(
        \i[20]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_19), .S(\i_4[20] ), .Y(), .FCO(i_4_cry_20));
    ARI1 #( .INIT(20'h42200) )  \i_RNIB7PP3[8]  (.A(VCC_net_1), .B(
        \i[8]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_7), .S(\i_4[8] ), .Y(), .FCO(i_4_cry_8));
    SLE \i[14]  (.D(\i_4[14] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[14]_net_1 ));
    SLE \i[0]  (.D(\i_4[0] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[0]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIA8TG4[19]  (.A(VCC_net_1), .B(
        \i[19]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_18), .S(\i_4[19] ), .Y(), .FCO(i_4_cry_19));
    SLE \i[13]  (.D(\i_4[13] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[13]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIK3OB4[15]  (.A(VCC_net_1), .B(
        \i[15]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_14), .S(\i_4[15] ), .Y(), .FCO(i_4_cry_15));
    CFG4 #( .INIT(16'h0008) )  un9_clklto22_i_0_a3 (.A(
        un9_clklto22_i_0_a3_1_net_1), .B(un9_clklto22_i_0_o2_net_1), 
        .C(\i[21]_net_1 ), .D(\i[20]_net_1 ), .Y(
        un9_clklto22_i_0_a3_net_1));
    SLE \i[5]  (.D(\i_4[5] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[5]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIS1H62[3]  (.A(VCC_net_1), .B(
        \i[3]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_2), .S(\i_4[3] ), .Y(), .FCO(i_4_cry_3));
    ARI1 #( .INIT(20'h42200) )  \i_RNI9GHJ4[21]  (.A(VCC_net_1), .B(
        \i[21]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_20), .S(\i_4[21] ), .Y(), .FCO(i_4_cry_21));
    ARI1 #( .INIT(20'h42200) )  \i_RNIT0PG2[4]  (.A(VCC_net_1), .B(
        \i[4]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_3), .S(\i_4[4] ), .Y(), .FCO(i_4_cry_4));
    SLE \i[16]  (.D(\i_4[16] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[16]_net_1 ));
    CFG4 #( .INIT(16'h7F77) )  un9_clklto22_i_0_o2_1 (.A(\i[9]_net_1 ), 
        .B(\i[8]_net_1 ), .C(\i[7]_net_1 ), .D(N_122), .Y(N_123));
    CFG4 #( .INIT(16'h5755) )  un9_clklto22_i_0_o2 (.A(\i[14]_net_1 ), 
        .B(\i[13]_net_1 ), .C(\i[12]_net_1 ), .D(N_124), .Y(
        un9_clklto22_i_0_o2_net_1));
    SLE \i[6]  (.D(\i_4[6] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[6]_net_1 ));
    SLE \i[19]  (.D(\i_4[19] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[19]_net_1 ));
    SLE \i[12]  (.D(\i_4[12] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[12]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \i_RNIJTJF4[18]  (.A(VCC_net_1), .B(
        \i[18]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_17), .S(\i_4[18] ), .Y(), .FCO(i_4_cry_18));
    CFG4 #( .INIT(16'h0007) )  un9_clklto22_i_0_a3_0 (.A(\i[19]_net_1 )
        , .B(\i[18]_net_1 ), .C(\i[21]_net_1 ), .D(\i[20]_net_1 ), .Y(
        un9_clklto22_i_0_a3_0_net_1));
    SLE \i[15]  (.D(\i_4[15] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[15]_net_1 ));
    ARI1 #( .INIT(20'h55500) )  \i_RNIVCA54[10]  (.A(\i[10]_net_1 ), 
        .B(pulse_meash_0_new_ready), .C(GND_net_1), .D(GND_net_1), 
        .FCI(i_4_cry_9), .S(\i_4[10] ), .Y(), .FCO(i_4_cry_10));
    CFG4 #( .INIT(16'h0F4F) )  un9_clklto22_i_0_o2_2 (.A(\i[0]_net_1 ), 
        .B(un9_clklto22_i_0_a2_2_3_net_1), .C(\i[6]_net_1 ), .D(
        \i[1]_net_1 ), .Y(N_122));
    ARI1 #( .INIT(20'h42200) )  \i_RNIV01R2[5]  (.A(VCC_net_1), .B(
        \i[5]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_4), .S(\i_4[5] ), .Y(), .FCO(i_4_cry_5));
    ARI1 #( .INIT(20'h42200) )  \i_RNI1TEA4[14]  (.A(VCC_net_1), .B(
        \i[14]_net_1 ), .C(pulse_meash_0_new_ready), .D(GND_net_1), 
        .FCI(i_4_cry_13), .S(\i_4[14] ), .Y(), .FCO(i_4_cry_14));
    SLE \i[7]  (.D(\i_4[7] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[7]_net_1 ));
    SLE \i[22]  (.D(\i_4[22] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[22]_net_1 ));
    SLE \i[4]  (.D(\i_4[4] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[4]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un9_clklto22_i_0_a2_2_3 (.A(
        \i[5]_net_1 ), .B(\i[4]_net_1 ), .C(\i[3]_net_1 ), .D(
        \i[2]_net_1 ), .Y(un9_clklto22_i_0_a2_2_3_net_1));
    SLE \i[1]  (.D(\i_4[1] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(\i[1]_net_1 ));
    SLE \i[11]  (.D(\i_4[11] ), .CLK(FCCC_0_GL0), .EN(FCCC_0_LOCK), 
        .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\i[11]_net_1 ));
    
endmodule


module Echo_control(
       LED_3_c,
       Echo_control_0_TX,
       mss_sb_0_TX,
       SERVO_PWM_c,
       ECHO_c,
       TRIG_c,
       LED_2_c
    );
output LED_3_c;
output Echo_control_0_TX;
input  mss_sb_0_TX;
output SERVO_PWM_c;
input  ECHO_c;
output TRIG_c;
output LED_2_c;

    wire \BT_module_0_data_buf[0] , \BT_module_0_data_buf[1] , 
        \BT_module_0_data_buf[2] , \BT_module_0_data_buf[3] , 
        \BT_module_0_data_buf[4] , \BT_module_0_data_buf[5] , 
        \BT_module_0_data_buf[6] , \BT_module_0_data_buf[7] , 
        \rx_dout_reg[0] , \rx_dout_reg[1] , \rx_dout_reg[2] , 
        \rx_dout_reg[3] , \rx_dout_reg[4] , \rx_dout_reg[5] , 
        \rx_dout_reg[6] , \rx_dout_reg[7] , FCCC_0_LOCK, FCCC_0_GL0, 
        BT_module_0_oen, COREUART_0_RXRDY, \time_sender_0_data_out[0] , 
        \time_sender_0_data_out[1] , \time_sender_0_data_out[2] , 
        \time_sender_0_data_out[3] , \time_sender_0_data_out[5] , 
        LED_3_c_i_0, COREUART_0_TXRDY, 
        OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC, 
        \locator_control_0_angle1[0] , \locator_control_0_angle1[1] , 
        \locator_control_0_angle1[2] , \locator_control_0_angle1[3] , 
        \pulse_meash_0_tim[0] , \pulse_meash_0_tim[1] , 
        \pulse_meash_0_tim[2] , \pulse_meash_0_tim[3] , 
        \pulse_meash_0_tim[4] , \pulse_meash_0_tim[5] , 
        \pulse_meash_0_tim[6] , \pulse_meash_0_tim[7] , 
        \pulse_meash_0_tim[8] , \pulse_meash_0_tim[9] , 
        \pulse_meash_0_tim[10] , \pulse_meash_0_tim[11] , 
        \pulse_meash_0_tim[12] , \pulse_meash_0_tim[13] , 
        pulse_meash_0_new_ready, un46_clk_0, un46_clk_1, un46_clk_2, 
        un46_clk_3, N_234_0, locator_control_0_en_timer, GND_net_1, 
        VCC_net_1;
    
    pulse_meash pulse_meash_0 (.pulse_meash_0_tim({
        \pulse_meash_0_tim[13] , \pulse_meash_0_tim[12] , 
        \pulse_meash_0_tim[11] , \pulse_meash_0_tim[10] , 
        \pulse_meash_0_tim[9] , \pulse_meash_0_tim[8] , 
        \pulse_meash_0_tim[7] , \pulse_meash_0_tim[6] , 
        \pulse_meash_0_tim[5] , \pulse_meash_0_tim[4] , 
        \pulse_meash_0_tim[3] , \pulse_meash_0_tim[2] , 
        \pulse_meash_0_tim[1] , \pulse_meash_0_tim[0] }), .FCCC_0_LOCK(
        FCCC_0_LOCK), .FCCC_0_GL0(FCCC_0_GL0), 
        .pulse_meash_0_new_ready(pulse_meash_0_new_ready), 
        .locator_control_0_en_timer(locator_control_0_en_timer), 
        .ECHO_c(ECHO_c));
    locator_control locator_control_0 (.BT_module_0_data_buf({
        \BT_module_0_data_buf[7] , \BT_module_0_data_buf[6] , 
        \BT_module_0_data_buf[5] , \BT_module_0_data_buf[4] , 
        \BT_module_0_data_buf[3] , \BT_module_0_data_buf[2] , 
        \BT_module_0_data_buf[1] , \BT_module_0_data_buf[0] }), 
        .locator_control_0_angle1({\locator_control_0_angle1[3] , 
        \locator_control_0_angle1[2] , \locator_control_0_angle1[1] , 
        \locator_control_0_angle1[0] }), .FCCC_0_LOCK(FCCC_0_LOCK), 
        .FCCC_0_GL0(FCCC_0_GL0), .un46_clk_0(un46_clk_0), .un46_clk_1(
        un46_clk_1), .un46_clk_2(un46_clk_2), .un46_clk_3(un46_clk_3), 
        .TRIG_c(TRIG_c), .locator_control_0_en_timer(
        locator_control_0_en_timer), .pulse_meash_0_new_ready(
        pulse_meash_0_new_ready), .N_234_0(N_234_0));
    time_sender time_sender_0 (.locator_control_0_angle1({
        \locator_control_0_angle1[3] , \locator_control_0_angle1[2] , 
        \locator_control_0_angle1[1] , \locator_control_0_angle1[0] }), 
        .pulse_meash_0_tim({\pulse_meash_0_tim[13] , 
        \pulse_meash_0_tim[12] , \pulse_meash_0_tim[11] , 
        \pulse_meash_0_tim[10] , \pulse_meash_0_tim[9] , 
        \pulse_meash_0_tim[8] , \pulse_meash_0_tim[7] , 
        \pulse_meash_0_tim[6] , \pulse_meash_0_tim[5] , 
        \pulse_meash_0_tim[4] , \pulse_meash_0_tim[3] , 
        \pulse_meash_0_tim[2] , \pulse_meash_0_tim[1] , 
        \pulse_meash_0_tim[0] }), .time_sender_0_data_out_0(
        \time_sender_0_data_out[0] ), .time_sender_0_data_out_1(
        \time_sender_0_data_out[1] ), .time_sender_0_data_out_2(
        \time_sender_0_data_out[2] ), .time_sender_0_data_out_3(
        \time_sender_0_data_out[3] ), .time_sender_0_data_out_5(
        \time_sender_0_data_out[5] ), .LED_3_c(LED_3_c), .LED_3_c_i_0(
        LED_3_c_i_0), .FCCC_0_GL0(FCCC_0_GL0), .FCCC_0_LOCK(
        FCCC_0_LOCK), .pulse_meash_0_new_ready(pulse_meash_0_new_ready)
        , .COREUART_0_TXRDY(COREUART_0_TXRDY));
    GND GND (.Y(GND_net_1));
    BT_module BT_module_0 (.BT_module_0_data_buf({
        \BT_module_0_data_buf[7] , \BT_module_0_data_buf[6] , 
        \BT_module_0_data_buf[5] , \BT_module_0_data_buf[4] , 
        \BT_module_0_data_buf[3] , \BT_module_0_data_buf[2] , 
        \BT_module_0_data_buf[1] , \BT_module_0_data_buf[0] }), 
        .rx_dout_reg({\rx_dout_reg[7] , \rx_dout_reg[6] , 
        \rx_dout_reg[5] , \rx_dout_reg[4] , \rx_dout_reg[3] , 
        \rx_dout_reg[2] , \rx_dout_reg[1] , \rx_dout_reg[0] }), 
        .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(FCCC_0_GL0), 
        .BT_module_0_oen(BT_module_0_oen), .COREUART_0_RXRDY(
        COREUART_0_RXRDY));
    servo_driver servo_driver_0 (.FCCC_0_LOCK(FCCC_0_LOCK), 
        .FCCC_0_GL0(FCCC_0_GL0), .SERVO_PWM_c(SERVO_PWM_c), 
        .un46_clk_0(un46_clk_0), .un46_clk_1(un46_clk_1), .un46_clk_2(
        un46_clk_2), .un46_clk_3(un46_clk_3), .N_234_0(N_234_0));
    VCC VCC (.Y(VCC_net_1));
    Echo_control_COREUART_0_COREUART_1s_1s_0s_19s_0s_0s COREUART_0 (
        .rx_dout_reg({\rx_dout_reg[7] , \rx_dout_reg[6] , 
        \rx_dout_reg[5] , \rx_dout_reg[4] , \rx_dout_reg[3] , 
        \rx_dout_reg[2] , \rx_dout_reg[1] , \rx_dout_reg[0] }), 
        .time_sender_0_data_out_0(\time_sender_0_data_out[0] ), 
        .time_sender_0_data_out_1(\time_sender_0_data_out[1] ), 
        .time_sender_0_data_out_2(\time_sender_0_data_out[2] ), 
        .time_sender_0_data_out_3(\time_sender_0_data_out[3] ), 
        .time_sender_0_data_out_5(\time_sender_0_data_out[5] ), 
        .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL0(FCCC_0_GL0), 
        .LED_3_c_i_0(LED_3_c_i_0), .COREUART_0_RXRDY(COREUART_0_RXRDY), 
        .LED_3_c(LED_3_c), .BT_module_0_oen(BT_module_0_oen), 
        .Echo_control_0_TX(Echo_control_0_TX), .COREUART_0_TXRDY(
        COREUART_0_TXRDY), .mss_sb_0_TX(mss_sb_0_TX));
    Echo_control_FCCC_0_FCCC FCCC_0 (.FCCC_0_LOCK(FCCC_0_LOCK), 
        .FCCC_0_GL0(FCCC_0_GL0), 
        .OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC(
        OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC));
    Echo_control_OSC_0_OSC OSC_0 (
        .OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC(
        OSC_0_RCOSC_1MHZ_CCC_OUT_RCOSC_1MHZ_CCC));
    delayer delayer_0 (.FCCC_0_GL0(FCCC_0_GL0), .FCCC_0_LOCK(
        FCCC_0_LOCK), .LED_2_c(LED_2_c), .pulse_meash_0_new_ready(
        pulse_meash_0_new_ready));
    
endmodule


module mss(
       PWM,
       BT_TX,
       DEVRST_N,
       ECHO,
       GPS_TX,
       BT_RX,
       GPS_RX,
       LED_1,
       LED_2,
       LED_3,
       SERVO_PWM,
       TRIG,
       COREI2C_0_0_SCL_IO,
       COREI2C_0_0_SDA_IO
    );
output [8:1] PWM;
input  BT_TX;
input  DEVRST_N;
input  ECHO;
input  GPS_TX;
output BT_RX;
output GPS_RX;
output LED_1;
output LED_2;
output LED_3;
output SERVO_PWM;
output TRIG;
inout  COREI2C_0_0_SCL_IO;
inout  COREI2C_0_0_SDA_IO;

    wire mss_sb_0_TX, Echo_control_0_TX, VCC_net_1, GND_net_1, BT_TX_c, 
        ECHO_c, GPS_TX_c, BT_RX_c, GPS_RX_c, LED_2_c, LED_3_c, 
        \PWM_c[1] , \PWM_c[2] , \PWM_c[3] , \PWM_c[4] , \PWM_c[5] , 
        \PWM_c[6] , \PWM_c[7] , \PWM_c[8] , SERVO_PWM_c, TRIG_c;
    
    OUTBUF BT_RX_obuf (.D(BT_RX_c), .PAD(BT_RX));
    OUTBUF \PWM_obuf[3]  (.D(\PWM_c[3] ), .PAD(PWM[3]));
    OUTBUF LED_1_obuf (.D(ECHO_c), .PAD(LED_1));
    mss_sb mss_sb_0 (.PWM_c({\PWM_c[8] , \PWM_c[7] , \PWM_c[6] , 
        \PWM_c[5] , \PWM_c[4] , \PWM_c[3] , \PWM_c[2] , \PWM_c[1] }), 
        .COREI2C_0_0_SDA_IO(COREI2C_0_0_SDA_IO), .COREI2C_0_0_SCL_IO(
        COREI2C_0_0_SCL_IO), .DEVRST_N(DEVRST_N), .mss_sb_0_TX(
        mss_sb_0_TX), .Echo_control_0_TX(Echo_control_0_TX), .GPS_RX_c(
        GPS_RX_c), .GPS_TX_c(GPS_TX_c), .BT_RX_c(BT_RX_c), .BT_TX_c(
        BT_TX_c));
    GND GND (.Y(GND_net_1));
    INBUF ECHO_ibuf (.PAD(ECHO), .Y(ECHO_c));
    OUTBUF \PWM_obuf[7]  (.D(\PWM_c[7] ), .PAD(PWM[7]));
    OUTBUF GPS_RX_obuf (.D(GPS_RX_c), .PAD(GPS_RX));
    Echo_control Echo_control_0 (.LED_3_c(LED_3_c), .Echo_control_0_TX(
        Echo_control_0_TX), .mss_sb_0_TX(mss_sb_0_TX), .SERVO_PWM_c(
        SERVO_PWM_c), .ECHO_c(ECHO_c), .TRIG_c(TRIG_c), .LED_2_c(
        LED_2_c));
    OUTBUF \PWM_obuf[1]  (.D(\PWM_c[1] ), .PAD(PWM[1]));
    OUTBUF \PWM_obuf[2]  (.D(\PWM_c[2] ), .PAD(PWM[2]));
    INBUF BT_TX_ibuf (.PAD(BT_TX), .Y(BT_TX_c));
    OUTBUF \PWM_obuf[6]  (.D(\PWM_c[6] ), .PAD(PWM[6]));
    OUTBUF \PWM_obuf[8]  (.D(\PWM_c[8] ), .PAD(PWM[8]));
    INBUF GPS_TX_ibuf (.PAD(GPS_TX), .Y(GPS_TX_c));
    OUTBUF SERVO_PWM_obuf (.D(SERVO_PWM_c), .PAD(SERVO_PWM));
    OUTBUF LED_3_obuf (.D(LED_3_c), .PAD(LED_3));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF \PWM_obuf[4]  (.D(\PWM_c[4] ), .PAD(PWM[4]));
    OUTBUF \PWM_obuf[5]  (.D(\PWM_c[5] ), .PAD(PWM[5]));
    OUTBUF TRIG_obuf (.D(TRIG_c), .PAD(TRIG));
    OUTBUF LED_2_obuf (.D(LED_2_c), .PAD(LED_2));
    
endmodule
